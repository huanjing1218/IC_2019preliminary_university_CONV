
module CONV_DW01_dec_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  CLKINVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  CLKINVX1 U2 ( .A(A[9]), .Y(n2) );
  OAI21XL U3 ( .A0(n3), .A1(n2), .B0(n4), .Y(SUM[9]) );
  AO21X1 U4 ( .A0(n5), .A1(A[8]), .B0(n3), .Y(SUM[8]) );
  OAI2BB1X1 U5 ( .A0N(n6), .A1N(A[7]), .B0(n5), .Y(SUM[7]) );
  OAI2BB1X1 U6 ( .A0N(n7), .A1N(A[6]), .B0(n6), .Y(SUM[6]) );
  OAI2BB1X1 U7 ( .A0N(n8), .A1N(A[5]), .B0(n7), .Y(SUM[5]) );
  OAI2BB1X1 U8 ( .A0N(n9), .A1N(A[4]), .B0(n8), .Y(SUM[4]) );
  OAI2BB1X1 U9 ( .A0N(n10), .A1N(A[3]), .B0(n9), .Y(SUM[3]) );
  OAI2BB1X1 U10 ( .A0N(n11), .A1N(A[2]), .B0(n10), .Y(SUM[2]) );
  OAI2BB1X1 U11 ( .A0N(A[0]), .A1N(A[1]), .B0(n11), .Y(SUM[1]) );
  XOR2X1 U12 ( .A(A[11]), .B(n12), .Y(SUM[11]) );
  NOR2X1 U13 ( .A(A[10]), .B(n4), .Y(n12) );
  XNOR2X1 U14 ( .A(A[10]), .B(n4), .Y(SUM[10]) );
  NAND2X1 U15 ( .A(n3), .B(n2), .Y(n4) );
  NOR2X1 U16 ( .A(n5), .B(A[8]), .Y(n3) );
  OR2X1 U17 ( .A(n6), .B(A[7]), .Y(n5) );
  OR2X1 U18 ( .A(n7), .B(A[6]), .Y(n6) );
  OR2X1 U19 ( .A(n8), .B(A[5]), .Y(n7) );
  OR2X1 U20 ( .A(n9), .B(A[4]), .Y(n8) );
  OR2X1 U21 ( .A(n10), .B(A[3]), .Y(n9) );
  OR2X1 U22 ( .A(n11), .B(A[2]), .Y(n10) );
  NAND2BX1 U23 ( .AN(A[1]), .B(SUM[0]), .Y(n11) );
endmodule


module CONV_DW_cmp_4 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [19:0] A;
  input [19:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181;

  NOR2BX1 U55 ( .AN(B[7]), .B(A[7]), .Y(n164) );
  OAI222X1 U56 ( .A0(B[5]), .A1(n130), .B0(B[5]), .B1(n169), .C0(n130), .C1(
        n169), .Y(n168) );
  CLKINVX1 U57 ( .A(A[12]), .Y(n126) );
  OAI222X1 U58 ( .A0(B[17]), .A1(n124), .B0(B[17]), .B1(n181), .C0(n181), .C1(
        n124), .Y(n180) );
  NAND2X1 U59 ( .A(n120), .B(n155), .Y(n149) );
  OA22X1 U60 ( .A0(B[10]), .A1(n127), .B0(B[10]), .B1(n161), .Y(n119) );
  AOI2BB2X2 U61 ( .B0(n143), .B1(n144), .A0N(n141), .A1N(n123), .Y(n142) );
  OAI222X1 U62 ( .A0(A[18]), .A1(n180), .B0(n180), .B1(n133), .C0(A[18]), .C1(
        n133), .Y(n141) );
  OAI21X1 U63 ( .A0(A[9]), .A1(n137), .B0(n163), .Y(n162) );
  NOR2BX1 U64 ( .AN(B[2]), .B(A[2]), .Y(n176) );
  OAI221X2 U65 ( .A0(B[19]), .A1(n141), .B0(B[19]), .B1(n123), .C0(n142), .Y(
        GE_LT_GT_LE) );
  NAND2BXL U66 ( .AN(B[7]), .B(A[7]), .Y(n179) );
  NAND2BXL U67 ( .AN(B[16]), .B(A[16]), .Y(n181) );
  NOR2BXL U68 ( .AN(B[16]), .B(A[16]), .Y(n147) );
  NAND2BXL U69 ( .AN(B[2]), .B(A[2]), .Y(n175) );
  AOI2BB1XL U70 ( .A0N(n140), .A1N(A[1]), .B0(B[0]), .Y(n177) );
  INVX1 U71 ( .A(B[18]), .Y(n133) );
  OAI222X4 U72 ( .A0(B[12]), .A1(n126), .B0(B[12]), .B1(n158), .C0(n158), .C1(
        n126), .Y(n157) );
  OAI222X4 U73 ( .A0(B[12]), .A1(n126), .B0(B[12]), .B1(n154), .C0(n126), .C1(
        n154), .Y(n153) );
  OR2X1 U74 ( .A(A[15]), .B(n134), .Y(n120) );
  NAND2X1 U75 ( .A(A[10]), .B(n128), .Y(n121) );
  NAND2X1 U76 ( .A(n159), .B(n160), .Y(n122) );
  AND3X2 U77 ( .A(n121), .B(n122), .C(n119), .Y(n148) );
  OAI21X4 U78 ( .A0(n148), .A1(n149), .B0(n150), .Y(n143) );
  OAI222X1 U79 ( .A0(A[15]), .A1(n151), .B0(n134), .B1(n151), .C0(A[15]), .C1(
        n134), .Y(n150) );
  OAI222X4 U80 ( .A0(B[14]), .A1(n125), .B0(B[14]), .B1(n152), .C0(n125), .C1(
        n152), .Y(n151) );
  CLKINVX1 U81 ( .A(A[5]), .Y(n130) );
  CLKINVX1 U82 ( .A(A[8]), .Y(n129) );
  CLKINVX1 U83 ( .A(A[17]), .Y(n124) );
  INVXL U84 ( .A(n175), .Y(n132) );
  OAI222X4 U85 ( .A0(A[13]), .A1(n157), .B0(n157), .B1(n135), .C0(A[13]), .C1(
        n135), .Y(n156) );
  OAI222X1 U86 ( .A0(A[9]), .A1(n178), .B0(n178), .B1(n137), .C0(A[9]), .C1(
        n137), .Y(n161) );
  INVX1 U87 ( .A(A[14]), .Y(n125) );
  OAI222X1 U88 ( .A0(A[13]), .A1(n153), .B0(n135), .B1(n153), .C0(A[13]), .C1(
        n135), .Y(n152) );
  NAND2X2 U89 ( .A(A[11]), .B(n136), .Y(n154) );
  OAI22XL U90 ( .A0(n156), .A1(n125), .B0(B[14]), .B1(n156), .Y(n155) );
  INVXL U91 ( .A(B[1]), .Y(n140) );
  CLKINVX1 U92 ( .A(A[3]), .Y(n131) );
  CLKINVX1 U93 ( .A(A[19]), .Y(n123) );
  CLKINVX1 U94 ( .A(A[10]), .Y(n127) );
  INVXL U95 ( .A(B[11]), .Y(n136) );
  INVXL U96 ( .A(B[4]), .Y(n139) );
  INVX1 U97 ( .A(B[13]), .Y(n135) );
  INVXL U98 ( .A(B[9]), .Y(n137) );
  INVXL U99 ( .A(B[6]), .Y(n138) );
  INVXL U100 ( .A(B[15]), .Y(n134) );
  OAI222X4 U101 ( .A0(B[8]), .A1(n129), .B0(B[8]), .B1(n179), .C0(n179), .C1(
        n129), .Y(n178) );
  INVX1 U102 ( .A(n161), .Y(n128) );
  OAI22XL U103 ( .A0(n123), .A1(n145), .B0(B[19]), .B1(n145), .Y(n144) );
  OAI21XL U104 ( .A0(A[18]), .A1(n133), .B0(n146), .Y(n145) );
  OAI22XL U105 ( .A0(n147), .A1(n124), .B0(B[17]), .B1(n147), .Y(n146) );
  NOR2X1 U106 ( .A(n136), .B(A[11]), .Y(n158) );
  OAI22XL U107 ( .A0(n127), .A1(n162), .B0(B[10]), .B1(n162), .Y(n160) );
  OAI22XL U108 ( .A0(n164), .A1(n129), .B0(B[8]), .B1(n164), .Y(n163) );
  OAI21XL U109 ( .A0(n165), .A1(n166), .B0(n167), .Y(n159) );
  OAI222XL U110 ( .A0(A[6]), .A1(n168), .B0(n138), .B1(n168), .C0(A[6]), .C1(
        n138), .Y(n167) );
  NAND2X1 U111 ( .A(A[4]), .B(n139), .Y(n169) );
  OAI21XL U112 ( .A0(A[6]), .A1(n138), .B0(n170), .Y(n166) );
  OAI22XL U113 ( .A0(n171), .A1(n130), .B0(B[5]), .B1(n171), .Y(n170) );
  NOR2X1 U114 ( .A(n139), .B(A[4]), .Y(n171) );
  AOI221XL U115 ( .A0(A[3]), .A1(n132), .B0(n172), .B1(n173), .C0(n174), .Y(
        n165) );
  OAI22XL U116 ( .A0(B[3]), .A1(n131), .B0(B[3]), .B1(n175), .Y(n174) );
  OAI22XL U117 ( .A0(n176), .A1(n131), .B0(B[3]), .B1(n176), .Y(n173) );
  AO22X1 U118 ( .A0(n177), .A1(A[0]), .B0(A[1]), .B1(n140), .Y(n172) );
endmodule


module CONV_DW01_inc_1 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2XL U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVXL U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module CONV_DW01_inc_2 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
endmodule


module CONV_DW_mult_tc_2 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n3, n5, n9, n12, n13, n15, n16, n17, n21, n22, n23, n24, n25, n27,
         n29, n30, n31, n33, n34, n35, n36, n40, n41, n43, n46, n47, n49, n51,
         n53, n54, n57, n58, n61, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n105, n106, n107, n108, n109, n111, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n130, n132, n134, n135, n136, n137, n138, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n174, n176, n179, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n203, n204, n205, n206,
         n207, n210, n211, n213, n215, n216, n218, n220, n221, n222, n223,
         n225, n227, n229, n232, n234, n235, n236, n237, n238, n240, n242,
         n244, n245, n246, n247, n248, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n309, n311, n312, n314, n315, n316,
         n318, n322, n323, n324, n325, n326, n332, n334, n335, n338, n339,
         n340, n341, n342, n343, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1044, n1046, n1049,
         n1050, n1058, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1091, n1092, n1094, n1098, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261;
  assign product[39] = n101;

  ADDFX2 U980 ( .A(n741), .B(n798), .CI(n623), .CO(n566), .S(n567) );
  OAI22X1 U981 ( .A0(n23), .A1(n971), .B0(n21), .B1(n970), .Y(n762) );
  NAND2X4 U982 ( .A(n1063), .B(n1083), .Y(n1073) );
  BUFX16 U983 ( .A(n1073), .Y(n41) );
  ADDFXL U984 ( .A(n372), .B(n646), .CI(n665), .CO(n365), .S(n366) );
  BUFX2 U985 ( .A(n1080), .Y(n58) );
  OA22XL U986 ( .A0(n1070), .A1(n845), .B0(n57), .B1(n844), .Y(n1225) );
  OAI22XL U987 ( .A0(n1070), .A1(n837), .B0(n58), .B1(n836), .Y(n372) );
  OR2X2 U988 ( .A(n1070), .B(n1215), .Y(n1211) );
  BUFX3 U989 ( .A(n765), .Y(n1186) );
  CLKBUFX3 U990 ( .A(n723), .Y(n1201) );
  OAI22X1 U991 ( .A0(n35), .A1(n932), .B0(n33), .B1(n931), .Y(n723) );
  BUFX2 U992 ( .A(n1087), .Y(n16) );
  OAI22X1 U993 ( .A0(n5), .A1(n1028), .B0(n1027), .B1(n3), .Y(n819) );
  BUFX6 U994 ( .A(n1089), .Y(n3) );
  OAI22X1 U995 ( .A0(n35), .A1(n933), .B0(n33), .B1(n932), .Y(n724) );
  OAI22X1 U996 ( .A0(n12), .A1(n1005), .B0(n9), .B1(n1004), .Y(n796) );
  BUFX6 U997 ( .A(n1088), .Y(n9) );
  XNOR2X2 U998 ( .A(n281), .B(n93), .Y(product[8]) );
  OAI22X1 U999 ( .A0(n17), .A1(n992), .B0(n15), .B1(n991), .Y(n783) );
  BUFX12 U1000 ( .A(n1077), .Y(n17) );
  CMPR42X2 U1001 ( .A(n779), .B(n1202), .C(n760), .D(n569), .ICI(n567), .S(
        n565), .ICO(n563), .CO(n564) );
  OAI22X1 U1002 ( .A0(n17), .A1(n988), .B0(n15), .B1(n987), .Y(n779) );
  CMPR42X2 U1003 ( .A(n725), .B(n763), .C(n801), .D(n820), .ICI(n595), .S(n591), .ICO(n589), .CO(n590) );
  OAI22X1 U1004 ( .A0(n23), .A1(n972), .B0(n21), .B1(n971), .Y(n763) );
  OAI22X1 U1005 ( .A0(n53), .A1(n870), .B0(n51), .B1(n869), .Y(n661) );
  BUFX4 U1006 ( .A(n1071), .Y(n53) );
  OAI21X2 U1007 ( .A0(n117), .A1(n115), .B0(n116), .Y(n114) );
  NOR2X2 U1008 ( .A(n1213), .B(n119), .Y(n117) );
  OAI22X1 U1009 ( .A0(n12), .A1(n1004), .B0(n9), .B1(n1003), .Y(n795) );
  BUFX20 U1010 ( .A(n1078), .Y(n12) );
  NAND2X2 U1011 ( .A(n1064), .B(n1084), .Y(n1074) );
  CLKBUFX3 U1012 ( .A(n1084), .Y(n33) );
  XNOR2X4 U1013 ( .A(a[9]), .B(a[10]), .Y(n1084) );
  BUFX8 U1014 ( .A(n49), .Y(n1183) );
  CLKBUFX2 U1015 ( .A(a[17]), .Y(n49) );
  OAI22X1 U1016 ( .A0(n47), .A1(n888), .B0(n46), .B1(n887), .Y(n679) );
  BUFX8 U1017 ( .A(n1072), .Y(n47) );
  ADDFHX2 U1018 ( .A(n704), .B(n742), .CI(n780), .CO(n576), .S(n577) );
  OAI22X1 U1019 ( .A0(n29), .A1(n951), .B0(n27), .B1(n950), .Y(n742) );
  CMPR42X2 U1020 ( .A(n696), .B(n658), .C(n810), .D(n1199), .ICI(n489), .S(
        n487), .ICO(n485), .CO(n486) );
  OAI22X1 U1021 ( .A0(n53), .A1(n867), .B0(n51), .B1(n866), .Y(n658) );
  ADDFX2 U1022 ( .A(n662), .B(n700), .CI(n757), .CO(n538), .S(n539) );
  ADDFHX2 U1023 ( .A(n718), .B(n794), .CI(n621), .CO(n525), .S(n526) );
  BUFX3 U1024 ( .A(n657), .Y(n1184) );
  OAI21X1 U1025 ( .A0(n109), .A1(n107), .B0(n108), .Y(n106) );
  AOI21X4 U1026 ( .A0(n114), .A1(n1196), .B0(n111), .Y(n109) );
  XNOR2XL U1027 ( .A(n734), .B(n639), .Y(n489) );
  OR2X2 U1028 ( .A(n734), .B(n639), .Y(n488) );
  OAI22X1 U1029 ( .A0(n1070), .A1(n848), .B0(n57), .B1(n847), .Y(n639) );
  INVX1 U1030 ( .A(n263), .Y(n262) );
  OAI21X4 U1031 ( .A0(n276), .A1(n264), .B0(n265), .Y(n263) );
  OAI22X1 U1032 ( .A0(n5), .A1(n1030), .B0(n1029), .B1(n3), .Y(n821) );
  BUFX20 U1033 ( .A(b[0]), .Y(n61) );
  OAI22X2 U1034 ( .A0(n5), .A1(n1238), .B0(n1039), .B1(n3), .Y(n629) );
  BUFX12 U1035 ( .A(n1079), .Y(n5) );
  BUFX6 U1036 ( .A(n404), .Y(n1185) );
  OAI22X1 U1037 ( .A0(n1070), .A1(n841), .B0(n57), .B1(n840), .Y(n404) );
  OAI22X4 U1038 ( .A0(n30), .A1(n1244), .B0(n27), .B1(n955), .Y(n625) );
  OAI22X1 U1039 ( .A0(n30), .A1(n943), .B0(n27), .B1(n942), .Y(n734) );
  OAI22X1 U1040 ( .A0(n30), .A1(n936), .B0(n27), .B1(n935), .Y(n727) );
  OAI22X1 U1041 ( .A0(n30), .A1(n942), .B0(n27), .B1(n941), .Y(n733) );
  CLKBUFX6 U1042 ( .A(n1075), .Y(n30) );
  BUFX4 U1043 ( .A(b[10]), .Y(n1049) );
  BUFX4 U1044 ( .A(b[15]), .Y(n1044) );
  INVX12 U1045 ( .A(n1232), .Y(n1233) );
  BUFX4 U1046 ( .A(b[19]), .Y(n1040) );
  XNOR2X1 U1047 ( .A(n1233), .B(b[2]), .Y(n994) );
  NOR2X2 U1048 ( .A(n194), .B(n191), .Y(n189) );
  CLKINVX3 U1049 ( .A(n292), .Y(n1236) );
  CLKAND2X8 U1050 ( .A(n1217), .B(n1200), .Y(n276) );
  AOI21X2 U1051 ( .A0(n186), .A1(n169), .B0(n170), .Y(n168) );
  OR2X1 U1052 ( .A(n542), .B(n552), .Y(n1191) );
  CLKINVX1 U1053 ( .A(n132), .Y(n130) );
  NAND2XL U1054 ( .A(n323), .B(n192), .Y(n78) );
  XNOR2X1 U1055 ( .A(n143), .B(n70), .Y(product[31]) );
  INVX3 U1056 ( .A(a[13]), .Y(n1209) );
  BUFX4 U1057 ( .A(a[15]), .Y(n43) );
  XOR2X1 U1058 ( .A(n620), .B(n792), .Y(n503) );
  OAI22XL U1059 ( .A0(n35), .A1(n927), .B0(n33), .B1(n926), .Y(n718) );
  OAI22XL U1060 ( .A0(n5), .A1(n1022), .B0(n1021), .B1(n3), .Y(n813) );
  OAI22XL U1061 ( .A0(n41), .A1(n909), .B0(n40), .B1(n908), .Y(n700) );
  INVX3 U1062 ( .A(n13), .Y(n1232) );
  INVX3 U1063 ( .A(n25), .Y(n1244) );
  CLKBUFX3 U1064 ( .A(b[13]), .Y(n1046) );
  CLKBUFX3 U1065 ( .A(n1080), .Y(n57) );
  CLKBUFX3 U1066 ( .A(b[18]), .Y(n1041) );
  OAI22XL U1067 ( .A0(n23), .A1(n967), .B0(n21), .B1(n966), .Y(n758) );
  OAI22XL U1068 ( .A0(n23), .A1(n975), .B0(n21), .B1(n974), .Y(n766) );
  NOR2X1 U1069 ( .A(n257), .B(n260), .Y(n255) );
  CLKBUFX3 U1070 ( .A(n722), .Y(n1202) );
  NAND2X1 U1071 ( .A(n134), .B(n1190), .Y(n127) );
  CMPR42X1 U1072 ( .A(n501), .B(n498), .C(n508), .D(n504), .ICI(n495), .S(n492), .ICO(n490), .CO(n491) );
  NAND2X1 U1073 ( .A(n1188), .B(n1192), .Y(n222) );
  OR2X1 U1074 ( .A(n1248), .B(n1249), .Y(n828) );
  XOR2X1 U1075 ( .A(n627), .B(n825), .Y(n615) );
  CMPR42X1 U1076 ( .A(n767), .B(n786), .C(n805), .D(n824), .ICI(n1198), .S(
        n611), .ICO(n609), .CO(n610) );
  CMPR42X1 U1077 ( .A(n802), .B(n598), .C(n602), .D(n596), .ICI(n599), .S(n594), .ICO(n592), .CO(n593) );
  CMPR42X1 U1078 ( .A(n743), .B(n624), .C(n589), .D(n590), .ICI(n583), .S(n580), .ICO(n578), .CO(n579) );
  OAI22XL U1079 ( .A0(n36), .A1(n1094), .B0(n34), .B1(n934), .Y(n624) );
  NOR2X1 U1080 ( .A(n165), .B(n160), .Y(n158) );
  NAND2X1 U1081 ( .A(n158), .B(n146), .Y(n144) );
  AOI21X1 U1082 ( .A0(n159), .A1(n146), .B0(n147), .Y(n145) );
  NOR2X1 U1083 ( .A(n438), .B(n428), .Y(n183) );
  NAND2X1 U1084 ( .A(n438), .B(n428), .Y(n184) );
  OAI21XL U1085 ( .A0(n124), .A1(n120), .B0(n121), .Y(n119) );
  OAI21XL U1086 ( .A0(n142), .A1(n136), .B0(n137), .Y(n135) );
  CLKINVX1 U1087 ( .A(n181), .Y(n179) );
  OR2X1 U1088 ( .A(n518), .B(n530), .Y(n1188) );
  OR2X1 U1089 ( .A(n531), .B(n541), .Y(n1192) );
  CLKINVX1 U1090 ( .A(n220), .Y(n218) );
  OR2X1 U1091 ( .A(n492), .B(n505), .Y(n1193) );
  OR2X2 U1092 ( .A(n427), .B(n417), .Y(n1189) );
  NOR2X1 U1093 ( .A(n376), .B(n381), .Y(n148) );
  NOR2X1 U1094 ( .A(n368), .B(n364), .Y(n136) );
  CLKBUFX3 U1095 ( .A(n829), .Y(n1203) );
  NAND2X1 U1096 ( .A(n1203), .B(n629), .Y(n307) );
  NOR2X2 U1097 ( .A(n1234), .B(n290), .Y(n288) );
  AND2X2 U1098 ( .A(n289), .B(n297), .Y(n1234) );
  OR2X2 U1099 ( .A(n1235), .B(n1236), .Y(n290) );
  CLKINVX1 U1100 ( .A(n274), .Y(n272) );
  OR2X1 U1101 ( .A(n588), .B(n593), .Y(n1194) );
  CLKINVX1 U1102 ( .A(n276), .Y(n275) );
  NOR2X1 U1103 ( .A(n580), .B(n587), .Y(n260) );
  XNOR2X1 U1104 ( .A(n1257), .B(n86), .Y(product[15]) );
  XOR2X1 U1105 ( .A(n109), .B(n64), .Y(product[37]) );
  XNOR2X1 U1106 ( .A(n1255), .B(n73), .Y(product[28]) );
  AO21X2 U1107 ( .A0(n167), .A1(n1214), .B0(n164), .Y(n1255) );
  XNOR2X1 U1108 ( .A(n1254), .B(n80), .Y(product[21]) );
  OAI21X1 U1109 ( .A0(n284), .A1(n282), .B0(n283), .Y(n281) );
  NAND2X1 U1110 ( .A(n338), .B(n1218), .Y(n1219) );
  CLKINVX1 U1111 ( .A(n279), .Y(n338) );
  OAI22X1 U1112 ( .A0(n17), .A1(n994), .B0(n15), .B1(n993), .Y(n785) );
  CLKBUFX3 U1113 ( .A(n766), .Y(n1187) );
  OAI22X1 U1114 ( .A0(n12), .A1(n1003), .B0(n9), .B1(n1002), .Y(n794) );
  OAI22X1 U1115 ( .A0(n1078), .A1(n1012), .B0(n9), .B1(n1011), .Y(n803) );
  OAI22X1 U1116 ( .A0(n12), .A1(n1009), .B0(n9), .B1(n1008), .Y(n800) );
  OAI22X1 U1117 ( .A0(n12), .A1(n1006), .B0(n9), .B1(n1005), .Y(n797) );
  OAI22X1 U1118 ( .A0(n12), .A1(n1010), .B0(n9), .B1(n1009), .Y(n801) );
  OAI22X1 U1119 ( .A0(n12), .A1(n1017), .B0(n9), .B1(n1016), .Y(n808) );
  OAI22X1 U1120 ( .A0(n5), .A1(n1032), .B0(n1031), .B1(n3), .Y(n823) );
  OAI22X1 U1121 ( .A0(n24), .A1(n1240), .B0(n22), .B1(n976), .Y(n626) );
  CLKBUFX3 U1122 ( .A(n1076), .Y(n24) );
  CMPR42X2 U1123 ( .A(n804), .B(n1187), .C(n785), .D(n608), .ICI(n609), .S(
        n606), .ICO(n604), .CO(n605) );
  OAI22X1 U1124 ( .A0(n1078), .A1(n1013), .B0(n9), .B1(n1012), .Y(n804) );
  OAI22X1 U1125 ( .A0(n5), .A1(n1031), .B0(n1030), .B1(n3), .Y(n822) );
  INVX12 U1126 ( .A(n1238), .Y(n1239) );
  INVX4 U1127 ( .A(a[1]), .Y(n1238) );
  NAND2X1 U1128 ( .A(n1062), .B(n1082), .Y(n1072) );
  OR2X1 U1129 ( .A(n359), .B(n363), .Y(n1190) );
  OR2X1 U1130 ( .A(n408), .B(n416), .Y(n1195) );
  INVX12 U1131 ( .A(n1244), .Y(n1245) );
  OR2X1 U1132 ( .A(n350), .B(n349), .Y(n1196) );
  OR2X1 U1133 ( .A(n630), .B(n346), .Y(n1197) );
  XNOR2X1 U1134 ( .A(a[15]), .B(a[16]), .Y(n1081) );
  BUFX4 U1135 ( .A(n1081), .Y(n51) );
  XNOR2X1 U1136 ( .A(a[13]), .B(a[14]), .Y(n1082) );
  INVX4 U1137 ( .A(n1215), .Y(n1216) );
  INVX3 U1138 ( .A(a[19]), .Y(n1215) );
  OR2X1 U1139 ( .A(n506), .B(n517), .Y(n1208) );
  AND2X2 U1140 ( .A(n627), .B(n825), .Y(n1198) );
  AND2X2 U1141 ( .A(n620), .B(n792), .Y(n1199) );
  NOR2X1 U1142 ( .A(n601), .B(n605), .Y(n279) );
  INVX8 U1143 ( .A(n1240), .Y(n1241) );
  INVX3 U1144 ( .A(a[7]), .Y(n1240) );
  INVX16 U1145 ( .A(n1209), .Y(n1210) );
  XNOR2X1 U1146 ( .A(a[7]), .B(a[8]), .Y(n1085) );
  BUFX4 U1147 ( .A(n1085), .Y(n27) );
  BUFX4 U1148 ( .A(n1083), .Y(n40) );
  NAND2X4 U1149 ( .A(n1228), .B(n1229), .Y(n1088) );
  AND2X2 U1150 ( .A(n1219), .B(n280), .Y(n1200) );
  CLKBUFX4 U1151 ( .A(n1237), .Y(n21) );
  NOR2X1 U1152 ( .A(n123), .B(n120), .Y(n118) );
  NAND2X1 U1153 ( .A(n169), .B(n125), .Y(n123) );
  XNOR2X1 U1154 ( .A(n1205), .B(n1050), .Y(n1008) );
  INVX16 U1155 ( .A(n1204), .Y(n1205) );
  CLKBUFX8 U1156 ( .A(a[11]), .Y(n31) );
  ADDHX1 U1157 ( .A(n661), .B(n813), .CO(n527), .S(n528) );
  BUFX2 U1158 ( .A(n1074), .Y(n36) );
  BUFX4 U1159 ( .A(n1075), .Y(n29) );
  CLKBUFX6 U1160 ( .A(n1074), .Y(n35) );
  ADDHX1 U1161 ( .A(n745), .B(n821), .CO(n597), .S(n598) );
  BUFX3 U1162 ( .A(n1087), .Y(n15) );
  XNOR2X2 U1163 ( .A(a[3]), .B(a[4]), .Y(n1087) );
  XOR2X1 U1164 ( .A(a[5]), .B(a[4]), .Y(n1067) );
  OAI22X1 U1165 ( .A0(n35), .A1(n930), .B0(n33), .B1(n929), .Y(n721) );
  OAI22X1 U1166 ( .A0(n23), .A1(n973), .B0(n21), .B1(n972), .Y(n764) );
  CLKBUFX4 U1167 ( .A(n1076), .Y(n23) );
  CMPR42X2 U1168 ( .A(n761), .B(n799), .C(n1201), .D(n818), .ICI(n577), .S(
        n575), .ICO(n573), .CO(n574) );
  OAI22X1 U1169 ( .A0(n23), .A1(n970), .B0(n21), .B1(n969), .Y(n761) );
  CLKINVX6 U1170 ( .A(a[3]), .Y(n1204) );
  OR2X1 U1171 ( .A(n12), .B(n1008), .Y(n1206) );
  OR2X1 U1172 ( .A(n9), .B(n1007), .Y(n1207) );
  NAND2X2 U1173 ( .A(n1206), .B(n1207), .Y(n799) );
  XNOR2XL U1174 ( .A(n1205), .B(n1049), .Y(n1007) );
  XOR2X1 U1175 ( .A(n185), .B(n77), .Y(product[24]) );
  CLKINVX1 U1176 ( .A(n186), .Y(n185) );
  XNOR2X4 U1177 ( .A(n1250), .B(n75), .Y(product[26]) );
  OR2XL U1178 ( .A(n58), .B(n850), .Y(n1212) );
  NAND2X1 U1179 ( .A(n1211), .B(n1212), .Y(n620) );
  OAI22X1 U1180 ( .A0(n12), .A1(n1001), .B0(n9), .B1(n1000), .Y(n792) );
  NAND2BXL U1181 ( .AN(n61), .B(n1216), .Y(n850) );
  OAI21X2 U1182 ( .A0(n196), .A1(n194), .B0(n195), .Y(n193) );
  NOR2X2 U1183 ( .A(n452), .B(n463), .Y(n194) );
  NAND2X2 U1184 ( .A(n1065), .B(n1085), .Y(n1075) );
  AND2X1 U1185 ( .A(n186), .B(n118), .Y(n1213) );
  XOR2X4 U1186 ( .A(n117), .B(n66), .Y(product[35]) );
  OR2XL U1187 ( .A(n398), .B(n407), .Y(n1214) );
  CMPR42X2 U1188 ( .A(n412), .B(n413), .C(n410), .D(n401), .ICI(n406), .S(n398), .ICO(n396), .CO(n397) );
  CMPR42X2 U1189 ( .A(n422), .B(n419), .C(n411), .D(n414), .ICI(n415), .S(n408), .ICO(n406), .CO(n407) );
  NAND2X2 U1190 ( .A(n285), .B(n277), .Y(n1217) );
  CLKINVX1 U1191 ( .A(n283), .Y(n1218) );
  NAND2X2 U1192 ( .A(n606), .B(n610), .Y(n283) );
  NAND2X1 U1193 ( .A(n601), .B(n605), .Y(n280) );
  OR2XL U1194 ( .A(n17), .B(n995), .Y(n1220) );
  OR2XL U1195 ( .A(n15), .B(n994), .Y(n1221) );
  NAND2X1 U1196 ( .A(n1220), .B(n1221), .Y(n786) );
  XNOR2X4 U1197 ( .A(a[11]), .B(a[12]), .Y(n1083) );
  AOI21X2 U1198 ( .A0(n143), .A1(n315), .B0(n140), .Y(n138) );
  NAND2X2 U1199 ( .A(n1243), .B(n145), .Y(n143) );
  OR2XL U1200 ( .A(n47), .B(n891), .Y(n1222) );
  OR2XL U1201 ( .A(n46), .B(n890), .Y(n1223) );
  NAND2X1 U1202 ( .A(n1222), .B(n1223), .Y(n682) );
  ADDHX2 U1203 ( .A(n682), .B(n815), .CO(n549), .S(n550) );
  XNOR2XL U1204 ( .A(n43), .B(n61), .Y(n891) );
  BUFX4 U1205 ( .A(n1082), .Y(n46) );
  OR2XL U1206 ( .A(n382), .B(n389), .Y(n1224) );
  CMPR42X2 U1207 ( .A(n649), .B(n391), .C(n392), .D(n385), .ICI(n388), .S(n382), .ICO(n380), .CO(n381) );
  CMPR42X2 U1208 ( .A(n399), .B(n395), .C(n400), .D(n393), .ICI(n396), .S(n390), .ICO(n388), .CO(n389) );
  NAND2X2 U1209 ( .A(n1061), .B(n1081), .Y(n1071) );
  XOR2X1 U1210 ( .A(a[15]), .B(a[14]), .Y(n1062) );
  NAND2X4 U1211 ( .A(n398), .B(n407), .Y(n166) );
  OAI21X2 U1212 ( .A0(n145), .A1(n127), .B0(n128), .Y(n126) );
  INVX1 U1213 ( .A(n254), .Y(n253) );
  INVX1 U1214 ( .A(n286), .Y(n340) );
  OAI21X2 U1215 ( .A0(n257), .A1(n261), .B0(n258), .Y(n256) );
  INVX3 U1216 ( .A(n256), .Y(n1231) );
  NOR2X1 U1217 ( .A(n291), .B(n295), .Y(n1235) );
  NAND2X1 U1218 ( .A(n617), .B(n618), .Y(n295) );
  XNOR2X2 U1219 ( .A(a[17]), .B(a[18]), .Y(n1080) );
  XOR2X4 U1220 ( .A(n1226), .B(n84), .Y(product[17]) );
  OA21X2 U1221 ( .A0(n235), .A1(n229), .B0(n234), .Y(n1226) );
  OAI22X1 U1222 ( .A0(n12), .A1(n1007), .B0(n9), .B1(n1006), .Y(n798) );
  NAND2X2 U1223 ( .A(a[1]), .B(a[2]), .Y(n1228) );
  NAND2X4 U1224 ( .A(n1238), .B(n1227), .Y(n1229) );
  CLKINVX2 U1225 ( .A(a[2]), .Y(n1227) );
  NAND2X4 U1226 ( .A(n1068), .B(n1088), .Y(n1078) );
  AOI21X1 U1227 ( .A0(n135), .A1(n1190), .B0(n130), .Y(n128) );
  XOR2X1 U1228 ( .A(n288), .B(n95), .Y(product[6]) );
  CLKAND2X12 U1229 ( .A(n1230), .B(n1231), .Y(n254) );
  NAND2X4 U1230 ( .A(n255), .B(n263), .Y(n1230) );
  CLKBUFX2 U1231 ( .A(a[5]), .Y(n13) );
  OAI2BB1XL U1232 ( .A0N(n106), .A1N(n1197), .B0(n105), .Y(n1261) );
  OAI21X4 U1233 ( .A0(n300), .A1(n298), .B0(n299), .Y(n297) );
  OAI21X4 U1234 ( .A0(n288), .A1(n286), .B0(n287), .Y(n285) );
  NOR2X4 U1235 ( .A(n613), .B(n616), .Y(n291) );
  NAND2X2 U1236 ( .A(n613), .B(n616), .Y(n292) );
  NAND2X2 U1237 ( .A(n1067), .B(n1087), .Y(n1077) );
  AO21X4 U1238 ( .A0(n182), .A1(n1189), .B0(n179), .Y(n1250) );
  NAND2X2 U1239 ( .A(n189), .B(n197), .Y(n187) );
  NOR2X1 U1240 ( .A(n291), .B(n294), .Y(n289) );
  NOR2X2 U1241 ( .A(n617), .B(n618), .Y(n294) );
  BUFX6 U1242 ( .A(n1086), .Y(n1237) );
  OR2XL U1243 ( .A(n185), .B(n183), .Y(n1247) );
  NAND2X2 U1244 ( .A(n1247), .B(n184), .Y(n182) );
  NOR2X1 U1245 ( .A(n398), .B(n407), .Y(n165) );
  XNOR2X4 U1246 ( .A(n1256), .B(n68), .Y(product[33]) );
  AO21XL U1247 ( .A0(n143), .A1(n134), .B0(n135), .Y(n1256) );
  NAND2X1 U1248 ( .A(n828), .B(n809), .Y(n304) );
  ADDFHX1 U1249 ( .A(n746), .B(n1186), .CI(n803), .CO(n602), .S(n603) );
  NAND2X2 U1250 ( .A(n1260), .B(n223), .Y(n221) );
  OR2XL U1251 ( .A(n168), .B(n144), .Y(n1243) );
  OA21X2 U1252 ( .A0(n210), .A1(n223), .B0(n211), .Y(n1253) );
  NAND2XL U1253 ( .A(n1189), .B(n181), .Y(n76) );
  XNOR2X1 U1254 ( .A(n182), .B(n76), .Y(product[25]) );
  OAI21X4 U1255 ( .A0(n237), .A1(n254), .B0(n238), .Y(n236) );
  INVXL U1256 ( .A(n141), .Y(n315) );
  NAND2X1 U1257 ( .A(n382), .B(n389), .Y(n154) );
  NOR2XL U1258 ( .A(n5), .B(n1037), .Y(n1248) );
  CLKBUFX2 U1259 ( .A(a[9]), .Y(n25) );
  AND2XL U1260 ( .A(n562), .B(n571), .Y(n1242) );
  CMPR42X2 U1261 ( .A(n573), .B(n576), .C(n574), .D(n570), .ICI(n565), .S(n562), .ICO(n560), .CO(n561) );
  CMPR42X2 U1262 ( .A(n584), .B(n581), .C(n578), .D(n582), .ICI(n575), .S(n572), .ICO(n570), .CO(n571) );
  OR2X2 U1263 ( .A(n210), .B(n222), .Y(n1252) );
  CLKINVX1 U1264 ( .A(n236), .Y(n235) );
  AO21XL U1265 ( .A0(n253), .A1(n244), .B0(n245), .Y(n1257) );
  INVXL U1266 ( .A(n136), .Y(n314) );
  NOR2X1 U1267 ( .A(n246), .B(n251), .Y(n244) );
  INVX1 U1268 ( .A(n1261), .Y(n101) );
  NAND2X1 U1269 ( .A(n369), .B(n375), .Y(n142) );
  NOR2X1 U1270 ( .A(n382), .B(n389), .Y(n153) );
  NAND2XL U1271 ( .A(n562), .B(n571), .Y(n252) );
  NAND2BXL U1272 ( .AN(n61), .B(n1239), .Y(n1039) );
  XNOR2X1 U1273 ( .A(n1239), .B(n1058), .Y(n1037) );
  XNOR2X1 U1274 ( .A(n1239), .B(b[2]), .Y(n1036) );
  OAI22X1 U1275 ( .A0(n5), .A1(n1024), .B0(n1023), .B1(n3), .Y(n815) );
  OAI22X1 U1276 ( .A0(n5), .A1(n1025), .B0(n1024), .B1(n3), .Y(n816) );
  OAI22X1 U1277 ( .A0(n5), .A1(n1027), .B0(n1026), .B1(n3), .Y(n818) );
  OR2XL U1278 ( .A(n246), .B(n252), .Y(n1246) );
  NAND2X1 U1279 ( .A(n1246), .B(n247), .Y(n245) );
  NOR2X4 U1280 ( .A(n553), .B(n561), .Y(n246) );
  NAND2X1 U1281 ( .A(n553), .B(n561), .Y(n247) );
  AOI21X2 U1282 ( .A0(n245), .A1(n1191), .B0(n240), .Y(n238) );
  NOR2X1 U1283 ( .A(n1036), .B(n3), .Y(n1249) );
  NOR2X1 U1284 ( .A(n828), .B(n809), .Y(n303) );
  INVXL U1285 ( .A(n236), .Y(n1251) );
  AOI21X1 U1286 ( .A0(n1193), .A1(n218), .B0(n213), .Y(n211) );
  OAI21X1 U1287 ( .A0(n160), .A1(n166), .B0(n161), .Y(n159) );
  OAI21X1 U1288 ( .A0(n191), .A1(n195), .B0(n192), .Y(n190) );
  INVXL U1289 ( .A(n1192), .Y(n229) );
  NAND2X1 U1290 ( .A(n1194), .B(n271), .Y(n264) );
  NAND2X1 U1291 ( .A(n439), .B(n451), .Y(n192) );
  INVXL U1292 ( .A(n257), .Y(n334) );
  INVXL U1293 ( .A(n260), .Y(n335) );
  NAND2X1 U1294 ( .A(n531), .B(n541), .Y(n234) );
  NAND2XL U1295 ( .A(n358), .B(n356), .Y(n121) );
  INVXL U1296 ( .A(n168), .Y(n167) );
  OAI21X1 U1297 ( .A0(n168), .A1(n156), .B0(n157), .Y(n155) );
  AOI21X4 U1298 ( .A0(n206), .A1(n197), .B0(n198), .Y(n196) );
  OAI21X4 U1299 ( .A0(n187), .A1(n207), .B0(n188), .Y(n186) );
  XNOR2X2 U1300 ( .A(n193), .B(n78), .Y(product[23]) );
  INVXL U1301 ( .A(n191), .Y(n323) );
  OA21X4 U1302 ( .A0(n1251), .A1(n1252), .B0(n1253), .Y(n207) );
  NAND2XL U1303 ( .A(n322), .B(n184), .Y(n77) );
  OAI21X2 U1304 ( .A0(n199), .A1(n205), .B0(n200), .Y(n198) );
  NOR2X2 U1305 ( .A(n199), .B(n204), .Y(n197) );
  AO21XL U1306 ( .A0(n206), .A1(n326), .B0(n203), .Y(n1254) );
  INVX1 U1307 ( .A(n215), .Y(n213) );
  NAND2XL U1308 ( .A(n1208), .B(n220), .Y(n83) );
  XNOR2X1 U1309 ( .A(n221), .B(n83), .Y(product[18]) );
  NAND2XL U1310 ( .A(n271), .B(n274), .Y(n92) );
  NAND2X2 U1311 ( .A(n478), .B(n491), .Y(n205) );
  NOR2X1 U1312 ( .A(n478), .B(n491), .Y(n204) );
  NAND2XL U1313 ( .A(n334), .B(n258), .Y(n89) );
  NOR2X1 U1314 ( .A(n594), .B(n600), .Y(n273) );
  CMPR42X2 U1315 ( .A(n523), .B(n512), .C(n520), .D(n516), .ICI(n509), .S(n506), .ICO(n504), .CO(n505) );
  NAND2XL U1316 ( .A(n335), .B(n261), .Y(n90) );
  NAND2XL U1317 ( .A(n340), .B(n287), .Y(n95) );
  CMPR42X2 U1318 ( .A(n461), .B(n465), .C(n466), .D(n455), .ICI(n462), .S(n452), .ICO(n450), .CO(n451) );
  CMPR42X2 U1319 ( .A(n470), .B(n473), .C(n480), .D(n476), .ICI(n467), .S(n464), .ICO(n462), .CO(n463) );
  NOR2X1 U1320 ( .A(n562), .B(n571), .Y(n251) );
  CMPR42X2 U1321 ( .A(n433), .B(n423), .C(n430), .D(n420), .ICI(n426), .S(n417), .ICO(n415), .CO(n416) );
  NOR2X1 U1322 ( .A(n369), .B(n375), .Y(n141) );
  NOR2X1 U1323 ( .A(n358), .B(n356), .Y(n120) );
  NOR2X1 U1324 ( .A(n355), .B(n351), .Y(n115) );
  NOR2X1 U1325 ( .A(n348), .B(n347), .Y(n107) );
  NOR2X1 U1326 ( .A(n572), .B(n579), .Y(n257) );
  NOR2X1 U1327 ( .A(n606), .B(n610), .Y(n282) );
  NOR2X1 U1328 ( .A(n619), .B(n827), .Y(n298) );
  OAI22X1 U1329 ( .A0(n1070), .A1(n847), .B0(n57), .B1(n846), .Y(n474) );
  NOR2X1 U1330 ( .A(n611), .B(n612), .Y(n286) );
  NAND2BXL U1331 ( .AN(n306), .B(n307), .Y(n100) );
  NOR2XL U1332 ( .A(n1203), .B(n629), .Y(n306) );
  AO21XL U1333 ( .A0(n24), .A1(n22), .B0(n956), .Y(n747) );
  AO21XL U1334 ( .A0(n36), .A1(n34), .B0(n914), .Y(n705) );
  AO21XL U1335 ( .A0(n47), .A1(n46), .B0(n872), .Y(n663) );
  ADDFXL U1336 ( .A(n643), .B(n353), .CI(n354), .CO(n350), .S(n351) );
  ADDFXL U1337 ( .A(n352), .B(n631), .CI(n642), .CO(n348), .S(n349) );
  AO21XL U1338 ( .A0(n54), .A1(n51), .B0(n851), .Y(n642) );
  OAI22X1 U1339 ( .A0(n1070), .A1(n831), .B0(n58), .B1(n830), .Y(n346) );
  AO21XL U1340 ( .A0(n1070), .A1(n58), .B0(n830), .Y(n630) );
  ADDHX1 U1341 ( .A(n703), .B(n817), .CO(n568), .S(n569) );
  OAI22X1 U1342 ( .A0(n5), .A1(n1026), .B0(n1025), .B1(n3), .Y(n817) );
  ADDHX1 U1343 ( .A(n626), .B(n823), .CO(n607), .S(n608) );
  ADDHX1 U1344 ( .A(n724), .B(n819), .CO(n584), .S(n585) );
  OAI22XL U1345 ( .A0(n5), .A1(n1038), .B0(n1037), .B1(n3), .Y(n829) );
  NOR2BXL U1346 ( .AN(n61), .B(n40), .Y(n704) );
  NOR2BXL U1347 ( .AN(n61), .B(n27), .Y(n746) );
  CMPR42X2 U1348 ( .A(n683), .B(n721), .C(n778), .D(n816), .ICI(n566), .S(n559), .ICO(n557), .CO(n558) );
  NOR2BXL U1349 ( .AN(n61), .B(n33), .Y(n725) );
  NOR2BXL U1350 ( .AN(n61), .B(n21), .Y(n767) );
  NOR2BXL U1351 ( .AN(n61), .B(n9), .Y(n809) );
  NOR2BXL U1352 ( .AN(n61), .B(n3), .Y(product[0]) );
  XNOR2X1 U1353 ( .A(a[5]), .B(a[6]), .Y(n1086) );
  NAND2X4 U1354 ( .A(n1066), .B(n1237), .Y(n1076) );
  CLKINVX1 U1355 ( .A(a[0]), .Y(n1089) );
  BUFX12 U1356 ( .A(b[1]), .Y(n1058) );
  BUFX12 U1357 ( .A(b[9]), .Y(n1050) );
  NAND2X4 U1358 ( .A(n1060), .B(n1080), .Y(n1070) );
  NOR2XL U1359 ( .A(n17), .B(n1232), .Y(n1258) );
  NOR2XL U1360 ( .A(n16), .B(n997), .Y(n1259) );
  OR2X1 U1361 ( .A(n1258), .B(n1259), .Y(n627) );
  OAI22X1 U1362 ( .A0(n5), .A1(n1034), .B0(n1033), .B1(n3), .Y(n825) );
  NAND2BXL U1363 ( .AN(n61), .B(n1233), .Y(n997) );
  OR2X4 U1364 ( .A(n235), .B(n222), .Y(n1260) );
  AOI21X2 U1365 ( .A0(n1188), .A1(n232), .B0(n225), .Y(n223) );
  CLKINVX1 U1366 ( .A(n159), .Y(n157) );
  CLKINVX1 U1367 ( .A(n158), .Y(n156) );
  NOR2X1 U1368 ( .A(n144), .B(n127), .Y(n125) );
  NAND2X1 U1369 ( .A(n1189), .B(n1195), .Y(n171) );
  CLKINVX1 U1370 ( .A(n207), .Y(n206) );
  NAND2X1 U1371 ( .A(n1188), .B(n227), .Y(n84) );
  XNOR2X1 U1372 ( .A(n206), .B(n81), .Y(product[20]) );
  NAND2X1 U1373 ( .A(n326), .B(n205), .Y(n81) );
  CLKINVX1 U1374 ( .A(n204), .Y(n326) );
  XNOR2X1 U1375 ( .A(n167), .B(n74), .Y(product[27]) );
  NAND2X1 U1376 ( .A(n1214), .B(n166), .Y(n74) );
  AOI21X1 U1377 ( .A0(n198), .A1(n189), .B0(n190), .Y(n188) );
  NAND2X1 U1378 ( .A(n1193), .B(n1208), .Y(n210) );
  OAI21X1 U1379 ( .A0(n171), .A1(n184), .B0(n172), .Y(n170) );
  AOI21X1 U1380 ( .A0(n179), .A1(n1195), .B0(n174), .Y(n172) );
  CLKINVX1 U1381 ( .A(n176), .Y(n174) );
  CLKINVX1 U1382 ( .A(n227), .Y(n225) );
  NAND2X1 U1383 ( .A(n318), .B(n161), .Y(n73) );
  CLKINVX1 U1384 ( .A(n160), .Y(n318) );
  NOR2X1 U1385 ( .A(n171), .B(n183), .Y(n169) );
  NAND2X1 U1386 ( .A(n325), .B(n200), .Y(n80) );
  CLKINVX1 U1387 ( .A(n199), .Y(n325) );
  NAND2X1 U1388 ( .A(n1195), .B(n176), .Y(n75) );
  XOR2X1 U1389 ( .A(n216), .B(n82), .Y(product[19]) );
  NAND2X1 U1390 ( .A(n1193), .B(n215), .Y(n82) );
  AOI21X1 U1391 ( .A0(n221), .A1(n1208), .B0(n218), .Y(n216) );
  CLKINVX1 U1392 ( .A(n183), .Y(n322) );
  XOR2X1 U1393 ( .A(n196), .B(n79), .Y(product[22]) );
  NAND2X1 U1394 ( .A(n324), .B(n195), .Y(n79) );
  CLKINVX1 U1395 ( .A(n194), .Y(n324) );
  CLKINVX1 U1396 ( .A(n205), .Y(n203) );
  CLKINVX1 U1397 ( .A(n166), .Y(n164) );
  XNOR2X1 U1398 ( .A(n253), .B(n88), .Y(product[13]) );
  NAND2X1 U1399 ( .A(n249), .B(n252), .Y(n88) );
  XNOR2X1 U1400 ( .A(n114), .B(n65), .Y(product[36]) );
  NAND2X1 U1401 ( .A(n1196), .B(n113), .Y(n65) );
  XNOR2X1 U1402 ( .A(n275), .B(n92), .Y(product[9]) );
  XNOR2X1 U1403 ( .A(n155), .B(n72), .Y(product[29]) );
  NAND2X1 U1404 ( .A(n1224), .B(n154), .Y(n72) );
  XNOR2X1 U1405 ( .A(n122), .B(n67), .Y(product[34]) );
  NAND2X1 U1406 ( .A(n312), .B(n121), .Y(n67) );
  OAI21XL U1407 ( .A0(n185), .A1(n123), .B0(n124), .Y(n122) );
  CLKINVX1 U1408 ( .A(n120), .Y(n312) );
  NAND2X1 U1409 ( .A(n315), .B(n142), .Y(n70) );
  XNOR2X1 U1410 ( .A(n106), .B(n63), .Y(product[38]) );
  NAND2X1 U1411 ( .A(n1197), .B(n105), .Y(n63) );
  AOI21X1 U1412 ( .A0(n1194), .A1(n272), .B0(n267), .Y(n265) );
  NOR2X2 U1413 ( .A(n464), .B(n477), .Y(n199) );
  NOR2X2 U1414 ( .A(n390), .B(n397), .Y(n160) );
  NOR2X2 U1415 ( .A(n439), .B(n451), .Y(n191) );
  CLKINVX1 U1416 ( .A(n113), .Y(n111) );
  OAI21XL U1417 ( .A0(n148), .A1(n154), .B0(n149), .Y(n147) );
  AOI21X1 U1418 ( .A0(n170), .A1(n125), .B0(n126), .Y(n124) );
  XOR2X1 U1419 ( .A(n138), .B(n69), .Y(product[32]) );
  NAND2X1 U1420 ( .A(n314), .B(n137), .Y(n69) );
  XOR2X1 U1421 ( .A(n150), .B(n71), .Y(product[30]) );
  NAND2X1 U1422 ( .A(n316), .B(n149), .Y(n71) );
  AOI21X1 U1423 ( .A0(n155), .A1(n1224), .B0(n152), .Y(n150) );
  CLKINVX1 U1424 ( .A(n148), .Y(n316) );
  NAND2X1 U1425 ( .A(n244), .B(n1191), .Y(n237) );
  NOR2X1 U1426 ( .A(n141), .B(n136), .Y(n134) );
  NOR2X1 U1427 ( .A(n148), .B(n153), .Y(n146) );
  NAND2X1 U1428 ( .A(n452), .B(n463), .Y(n195) );
  NAND2X1 U1429 ( .A(n506), .B(n517), .Y(n220) );
  NAND2X1 U1430 ( .A(n408), .B(n416), .Y(n176) );
  NAND2X1 U1431 ( .A(n518), .B(n530), .Y(n227) );
  NAND2X1 U1432 ( .A(n492), .B(n505), .Y(n215) );
  NAND2X1 U1433 ( .A(n427), .B(n417), .Y(n181) );
  NAND2X1 U1434 ( .A(n464), .B(n477), .Y(n200) );
  NAND2X1 U1435 ( .A(n390), .B(n397), .Y(n161) );
  XOR2X1 U1436 ( .A(n270), .B(n91), .Y(product[10]) );
  NAND2X1 U1437 ( .A(n1194), .B(n269), .Y(n91) );
  AOI21X1 U1438 ( .A0(n275), .A1(n271), .B0(n272), .Y(n270) );
  XOR2X1 U1439 ( .A(n248), .B(n87), .Y(product[14]) );
  NAND2X1 U1440 ( .A(n332), .B(n247), .Y(n87) );
  AOI21X1 U1441 ( .A0(n253), .A1(n249), .B0(n1242), .Y(n248) );
  CLKINVX1 U1442 ( .A(n246), .Y(n332) );
  NAND2X1 U1443 ( .A(n1191), .B(n242), .Y(n86) );
  XOR2X1 U1444 ( .A(n235), .B(n85), .Y(product[16]) );
  NAND2X1 U1445 ( .A(n1192), .B(n234), .Y(n85) );
  NAND2X1 U1446 ( .A(n1190), .B(n132), .Y(n68) );
  NAND2X1 U1447 ( .A(n309), .B(n108), .Y(n64) );
  CLKINVX1 U1448 ( .A(n107), .Y(n309) );
  NAND2X1 U1449 ( .A(n311), .B(n116), .Y(n66) );
  CLKINVX1 U1450 ( .A(n115), .Y(n311) );
  CLKINVX1 U1451 ( .A(n273), .Y(n271) );
  CLKINVX1 U1452 ( .A(n234), .Y(n232) );
  CLKINVX1 U1453 ( .A(n285), .Y(n284) );
  CLKINVX1 U1454 ( .A(n297), .Y(n296) );
  CLKINVX1 U1455 ( .A(n251), .Y(n249) );
  CLKINVX1 U1456 ( .A(n269), .Y(n267) );
  CLKINVX1 U1457 ( .A(n242), .Y(n240) );
  CLKINVX1 U1458 ( .A(n142), .Y(n140) );
  CLKINVX1 U1459 ( .A(n154), .Y(n152) );
  XNOR2X1 U1460 ( .A(n99), .B(n305), .Y(product[2]) );
  NAND2X1 U1461 ( .A(n301), .B(n304), .Y(n99) );
  CMPR42X1 U1462 ( .A(n547), .B(n544), .C(n537), .D(n534), .ICI(n540), .S(n531), .ICO(n529), .CO(n530) );
  CMPR42X1 U1463 ( .A(n445), .B(n453), .C(n454), .D(n442), .ICI(n450), .S(n439), .ICO(n437), .CO(n438) );
  CMPR42X1 U1464 ( .A(n444), .B(n434), .C(n431), .D(n441), .ICI(n437), .S(n428), .ICO(n426), .CO(n427) );
  NOR2X1 U1465 ( .A(n279), .B(n282), .Y(n277) );
  AOI21X1 U1466 ( .A0(n301), .A1(n305), .B0(n302), .Y(n300) );
  CLKINVX1 U1467 ( .A(n304), .Y(n302) );
  CLKINVX1 U1468 ( .A(n303), .Y(n301) );
  NAND2X1 U1469 ( .A(n338), .B(n280), .Y(n93) );
  XNOR2X1 U1470 ( .A(n259), .B(n89), .Y(product[12]) );
  OAI21XL U1471 ( .A0(n262), .A1(n260), .B0(n261), .Y(n259) );
  NAND2X1 U1472 ( .A(n542), .B(n552), .Y(n242) );
  NAND2X1 U1473 ( .A(n594), .B(n600), .Y(n274) );
  NAND2X1 U1474 ( .A(n588), .B(n593), .Y(n269) );
  NAND2X1 U1475 ( .A(n376), .B(n381), .Y(n149) );
  XOR2X1 U1476 ( .A(n98), .B(n300), .Y(product[3]) );
  NAND2X1 U1477 ( .A(n343), .B(n299), .Y(n98) );
  CLKINVX1 U1478 ( .A(n298), .Y(n343) );
  XOR2X1 U1479 ( .A(n262), .B(n90), .Y(product[11]) );
  XOR2X1 U1480 ( .A(n296), .B(n97), .Y(product[4]) );
  NAND2X1 U1481 ( .A(n342), .B(n295), .Y(n97) );
  CLKINVX1 U1482 ( .A(n294), .Y(n342) );
  XOR2X1 U1483 ( .A(n284), .B(n94), .Y(product[7]) );
  NAND2X1 U1484 ( .A(n339), .B(n283), .Y(n94) );
  CLKINVX1 U1485 ( .A(n282), .Y(n339) );
  CMPR42X1 U1486 ( .A(n536), .B(n533), .C(n524), .D(n521), .ICI(n529), .S(n518), .ICO(n516), .CO(n517) );
  CMPR42X1 U1487 ( .A(n484), .B(n487), .C(n494), .D(n490), .ICI(n481), .S(n478), .ICO(n476), .CO(n477) );
  CLKINVX1 U1488 ( .A(n307), .Y(n305) );
  CLKINVX1 U1489 ( .A(n474), .Y(n475) );
  XNOR2X1 U1490 ( .A(n293), .B(n96), .Y(product[5]) );
  OAI21XL U1491 ( .A0(n296), .A1(n294), .B0(n295), .Y(n293) );
  NAND2X1 U1492 ( .A(n341), .B(n292), .Y(n96) );
  CLKINVX1 U1493 ( .A(n291), .Y(n341) );
  NAND2X1 U1494 ( .A(n359), .B(n363), .Y(n132) );
  NAND2X1 U1495 ( .A(n368), .B(n364), .Y(n137) );
  NAND2X1 U1496 ( .A(n355), .B(n351), .Y(n116) );
  NAND2X1 U1497 ( .A(n350), .B(n349), .Y(n113) );
  CLKINVX1 U1498 ( .A(n346), .Y(n347) );
  NAND2X1 U1499 ( .A(n348), .B(n347), .Y(n108) );
  NAND2X1 U1500 ( .A(n630), .B(n346), .Y(n105) );
  OAI22XL U1501 ( .A0(n1070), .A1(n845), .B0(n57), .B1(n844), .Y(n448) );
  OAI22X1 U1502 ( .A0(n1070), .A1(n843), .B0(n57), .B1(n842), .Y(n424) );
  OAI22X1 U1503 ( .A0(n1070), .A1(n839), .B0(n58), .B1(n838), .Y(n386) );
  OAI22XL U1504 ( .A0(n5), .A1(n1036), .B0(n1035), .B1(n3), .Y(n827) );
  CMPR42X1 U1505 ( .A(n784), .B(n822), .C(n607), .D(n604), .ICI(n603), .S(n601), .ICO(n599), .CO(n600) );
  OAI22XL U1506 ( .A0(n17), .A1(n993), .B0(n15), .B1(n992), .Y(n784) );
  CMPR42X1 U1507 ( .A(n558), .B(n555), .C(n545), .D(n548), .ICI(n551), .S(n542), .ICO(n540), .CO(n541) );
  OAI22XL U1508 ( .A0(n54), .A1(n858), .B0(n51), .B1(n857), .Y(n649) );
  CMPR42X1 U1509 ( .A(n685), .B(n377), .C(n371), .D(n378), .ICI(n374), .S(n369), .ICO(n367), .CO(n368) );
  OAI22XL U1510 ( .A0(n1073), .A1(n894), .B0(n40), .B1(n893), .Y(n685) );
  CMPR42X1 U1511 ( .A(n634), .B(n648), .C(n384), .D(n379), .ICI(n380), .S(n376), .ICO(n374), .CO(n375) );
  OAI22XL U1512 ( .A0(n54), .A1(n857), .B0(n51), .B1(n856), .Y(n648) );
  OAI22XL U1513 ( .A0(n1070), .A1(n838), .B0(n58), .B1(n837), .Y(n634) );
  CMPR42X1 U1514 ( .A(n782), .B(n744), .C(n597), .D(n592), .ICI(n591), .S(n588), .ICO(n586), .CO(n587) );
  OAI22XL U1515 ( .A0(n29), .A1(n953), .B0(n27), .B1(n952), .Y(n744) );
  OAI22XL U1516 ( .A0(n17), .A1(n991), .B0(n15), .B1(n990), .Y(n782) );
  CMPR42X1 U1517 ( .A(n568), .B(n559), .C(n564), .D(n556), .ICI(n560), .S(n553), .ICO(n551), .CO(n552) );
  OAI22XL U1518 ( .A0(n36), .A1(n918), .B0(n34), .B1(n917), .Y(n709) );
  OAI22XL U1519 ( .A0(n41), .A1(n910), .B0(n40), .B1(n909), .Y(n701) );
  OAI22XL U1520 ( .A0(n41), .A1(n906), .B0(n1083), .B1(n905), .Y(n697) );
  OAI22XL U1521 ( .A0(n12), .A1(n1000), .B0(n9), .B1(n999), .Y(n791) );
  OAI22XL U1522 ( .A0(n41), .A1(n905), .B0(n1083), .B1(n904), .Y(n696) );
  OAI22XL U1523 ( .A0(n12), .A1(n1002), .B0(n9), .B1(n1001), .Y(n793) );
  OAI22XL U1524 ( .A0(n1070), .A1(n846), .B0(n57), .B1(n845), .Y(n638) );
  OAI22XL U1525 ( .A0(n1070), .A1(n844), .B0(n57), .B1(n843), .Y(n637) );
  OAI22XL U1526 ( .A0(n24), .A1(n959), .B0(n22), .B1(n958), .Y(n750) );
  OAI22XL U1527 ( .A0(n1073), .A1(n900), .B0(n40), .B1(n899), .Y(n691) );
  OAI22XL U1528 ( .A0(n47), .A1(n877), .B0(n46), .B1(n876), .Y(n668) );
  OAI22XL U1529 ( .A0(n1070), .A1(n840), .B0(n57), .B1(n839), .Y(n635) );
  CMPR42X1 U1530 ( .A(n708), .B(n651), .C(n689), .D(n409), .ICI(n403), .S(n401), .ICO(n399), .CO(n400) );
  OAI22XL U1531 ( .A0(n1073), .A1(n898), .B0(n40), .B1(n897), .Y(n689) );
  OAI22XL U1532 ( .A0(n54), .A1(n860), .B0(n51), .B1(n859), .Y(n651) );
  OAI22XL U1533 ( .A0(n36), .A1(n917), .B0(n34), .B1(n916), .Y(n708) );
  CLKINVX1 U1534 ( .A(n100), .Y(product[1]) );
  NAND2X1 U1535 ( .A(n580), .B(n587), .Y(n261) );
  CMPR42X1 U1536 ( .A(n697), .B(n754), .C(n659), .D(n678), .ICI(n510), .S(n498), .ICO(n496), .CO(n497) );
  OAI22XL U1537 ( .A0(n47), .A1(n887), .B0(n46), .B1(n886), .Y(n678) );
  OAI22XL U1538 ( .A0(n53), .A1(n868), .B0(n51), .B1(n867), .Y(n659) );
  OAI22XL U1539 ( .A0(n24), .A1(n963), .B0(n22), .B1(n962), .Y(n754) );
  CMPR42X1 U1540 ( .A(n793), .B(n660), .C(n774), .D(n736), .ICI(n522), .S(n512), .ICO(n510), .CO(n511) );
  OAI22XL U1541 ( .A0(n29), .A1(n945), .B0(n27), .B1(n944), .Y(n736) );
  OAI22XL U1542 ( .A0(n1077), .A1(n983), .B0(n16), .B1(n982), .Y(n774) );
  OAI22XL U1543 ( .A0(n53), .A1(n869), .B0(n51), .B1(n868), .Y(n660) );
  CMPR42X1 U1544 ( .A(n640), .B(n773), .C(n811), .D(n503), .ICI(n507), .S(n501), .ICO(n499), .CO(n500) );
  OAI22XL U1545 ( .A0(n5), .A1(n1020), .B0(n1019), .B1(n3), .Y(n811) );
  OAI22XL U1546 ( .A0(n17), .A1(n982), .B0(n16), .B1(n981), .Y(n773) );
  OAI22XL U1547 ( .A0(n1070), .A1(n849), .B0(n57), .B1(n848), .Y(n640) );
  CMPR42X1 U1548 ( .A(n750), .B(n655), .C(n731), .D(n674), .ICI(n447), .S(n445), .ICO(n443), .CO(n444) );
  OAI22XL U1549 ( .A0(n47), .A1(n883), .B0(n46), .B1(n882), .Y(n674) );
  OAI22XL U1550 ( .A0(n30), .A1(n940), .B0(n27), .B1(n939), .Y(n731) );
  OAI22XL U1551 ( .A0(n53), .A1(n864), .B0(n51), .B1(n863), .Y(n655) );
  CMPR42X1 U1552 ( .A(n719), .B(n681), .C(n549), .D(n543), .ICI(n546), .S(n534), .ICO(n532), .CO(n533) );
  OAI22XL U1553 ( .A0(n47), .A1(n890), .B0(n46), .B1(n889), .Y(n681) );
  OAI22XL U1554 ( .A0(n35), .A1(n928), .B0(n33), .B1(n927), .Y(n719) );
  CMPR42X1 U1555 ( .A(n424), .B(n728), .C(n671), .D(n747), .ICI(n421), .S(n414), .ICO(n412), .CO(n413) );
  OAI22XL U1556 ( .A0(n47), .A1(n880), .B0(n46), .B1(n879), .Y(n671) );
  OAI22XL U1557 ( .A0(n30), .A1(n937), .B0(n27), .B1(n936), .Y(n728) );
  CMPR42X1 U1558 ( .A(n729), .B(n672), .C(n710), .D(n432), .ICI(n429), .S(n420), .ICO(n418), .CO(n419) );
  OAI22XL U1559 ( .A0(n36), .A1(n919), .B0(n34), .B1(n918), .Y(n710) );
  OAI22XL U1560 ( .A0(n47), .A1(n881), .B0(n46), .B1(n880), .Y(n672) );
  OAI22XL U1561 ( .A0(n30), .A1(n938), .B0(n27), .B1(n937), .Y(n729) );
  CMPR42X1 U1562 ( .A(n739), .B(n796), .C(n777), .D(n550), .ICI(n554), .S(n548), .ICO(n546), .CO(n547) );
  OAI22XL U1563 ( .A0(n17), .A1(n986), .B0(n16), .B1(n985), .Y(n777) );
  OAI22XL U1564 ( .A0(n29), .A1(n948), .B0(n27), .B1(n947), .Y(n739) );
  CMPR42X1 U1565 ( .A(n637), .B(n673), .C(n730), .D(n768), .ICI(n446), .S(n434), .ICO(n432), .CO(n433) );
  AO21X1 U1566 ( .A0(n1077), .A1(n16), .B0(n977), .Y(n768) );
  OAI22XL U1567 ( .A0(n30), .A1(n939), .B0(n27), .B1(n938), .Y(n730) );
  OAI22XL U1568 ( .A0(n47), .A1(n882), .B0(n46), .B1(n881), .Y(n673) );
  CMPR42X1 U1569 ( .A(n691), .B(n748), .C(n653), .D(n425), .ICI(n435), .S(n423), .ICO(n421), .CO(n422) );
  OAI22XL U1570 ( .A0(n53), .A1(n862), .B0(n51), .B1(n861), .Y(n653) );
  CLKINVX1 U1571 ( .A(n424), .Y(n425) );
  OAI22XL U1572 ( .A0(n24), .A1(n957), .B0(n22), .B1(n956), .Y(n748) );
  CMPR42X1 U1573 ( .A(n711), .B(n692), .C(n443), .D(n436), .ICI(n440), .S(n431), .ICO(n429), .CO(n430) );
  OAI22XL U1574 ( .A0(n1073), .A1(n901), .B0(n40), .B1(n900), .Y(n692) );
  OAI22XL U1575 ( .A0(n36), .A1(n920), .B0(n34), .B1(n919), .Y(n711) );
  CMPR42X1 U1576 ( .A(n701), .B(n758), .C(n622), .D(n720), .ICI(n557), .S(n545), .ICO(n543), .CO(n544) );
  OAI22XL U1577 ( .A0(n35), .A1(n929), .B0(n33), .B1(n928), .Y(n720) );
  OAI22XL U1578 ( .A0(n47), .A1(n1092), .B0(n46), .B1(n892), .Y(n622) );
  CMPR42X1 U1579 ( .A(n775), .B(n680), .C(n699), .D(n528), .ICI(n532), .S(n524), .ICO(n522), .CO(n523) );
  OAI22XL U1580 ( .A0(n41), .A1(n908), .B0(n1083), .B1(n907), .Y(n699) );
  OAI22XL U1581 ( .A0(n47), .A1(n889), .B0(n46), .B1(n888), .Y(n680) );
  OAI22XL U1582 ( .A0(n17), .A1(n984), .B0(n16), .B1(n983), .Y(n775) );
  NAND2X1 U1583 ( .A(n611), .B(n612), .Y(n287) );
  NAND2X1 U1584 ( .A(n572), .B(n579), .Y(n258) );
  CMPR42X1 U1585 ( .A(n738), .B(n795), .C(n776), .D(n814), .ICI(n539), .S(n537), .ICO(n535), .CO(n536) );
  OAI22XL U1586 ( .A0(n5), .A1(n1023), .B0(n1022), .B1(n3), .Y(n814) );
  OAI22XL U1587 ( .A0(n17), .A1(n985), .B0(n16), .B1(n984), .Y(n776) );
  OAI22XL U1588 ( .A0(n29), .A1(n947), .B0(n27), .B1(n946), .Y(n738) );
  CMPR42X1 U1589 ( .A(n717), .B(n698), .C(n527), .D(n519), .ICI(n515), .S(n509), .ICO(n507), .CO(n508) );
  OAI22XL U1590 ( .A0(n41), .A1(n907), .B0(n1083), .B1(n906), .Y(n698) );
  OAI22XL U1591 ( .A0(n35), .A1(n926), .B0(n33), .B1(n925), .Y(n717) );
  CMPR42X1 U1592 ( .A(n695), .B(n1184), .C(n475), .D(n488), .ICI(n485), .S(
        n473), .ICO(n471), .CO(n472) );
  OAI22XL U1593 ( .A0(n53), .A1(n866), .B0(n51), .B1(n865), .Y(n657) );
  OAI22XL U1594 ( .A0(n41), .A1(n904), .B0(n40), .B1(n903), .Y(n695) );
  OAI22XL U1595 ( .A0(n23), .A1(n969), .B0(n21), .B1(n968), .Y(n760) );
  OAI22XL U1596 ( .A0(n35), .A1(n931), .B0(n33), .B1(n930), .Y(n722) );
  AO21X1 U1597 ( .A0(n1079), .A1(n3), .B0(n1019), .Y(n810) );
  CMPR42X1 U1598 ( .A(n737), .B(n756), .C(n535), .D(n538), .ICI(n526), .S(n521), .ICO(n519), .CO(n520) );
  OAI22XL U1599 ( .A0(n24), .A1(n965), .B0(n22), .B1(n964), .Y(n756) );
  OAI22XL U1600 ( .A0(n29), .A1(n946), .B0(n27), .B1(n945), .Y(n737) );
  CMPR42X1 U1601 ( .A(n753), .B(n499), .C(n493), .D(n500), .ICI(n497), .S(n481), .ICO(n479), .CO(n480) );
  OAI22XL U1602 ( .A0(n24), .A1(n962), .B0(n22), .B1(n961), .Y(n753) );
  CMPR42X1 U1603 ( .A(n714), .B(n676), .C(n486), .D(n483), .ICI(n479), .S(n467), .ICO(n465), .CO(n466) );
  OAI22XL U1604 ( .A0(n47), .A1(n885), .B0(n46), .B1(n884), .Y(n676) );
  OAI22XL U1605 ( .A0(n36), .A1(n923), .B0(n34), .B1(n922), .Y(n714) );
  CMPR42X1 U1606 ( .A(n668), .B(n706), .C(n687), .D(n387), .ICI(n394), .S(n385), .ICO(n383), .CO(n384) );
  OAI22XL U1607 ( .A0(n41), .A1(n896), .B0(n40), .B1(n895), .Y(n687) );
  OAI22XL U1608 ( .A0(n36), .A1(n915), .B0(n34), .B1(n914), .Y(n706) );
  CLKINVX1 U1609 ( .A(n386), .Y(n387) );
  CMPR42X1 U1610 ( .A(n635), .B(n688), .C(n669), .D(n726), .ICI(n402), .S(n393), .ICO(n391), .CO(n392) );
  AO21X1 U1611 ( .A0(n30), .A1(n27), .B0(n935), .Y(n726) );
  OAI22XL U1612 ( .A0(n47), .A1(n878), .B0(n46), .B1(n877), .Y(n669) );
  OAI22XL U1613 ( .A0(n1073), .A1(n897), .B0(n40), .B1(n896), .Y(n688) );
  CMPR42X1 U1614 ( .A(n386), .B(n686), .C(n667), .D(n705), .ICI(n383), .S(n379), .ICO(n377), .CO(n378) );
  OAI22XL U1615 ( .A0(n47), .A1(n876), .B0(n46), .B1(n875), .Y(n667) );
  OAI22XL U1616 ( .A0(n41), .A1(n895), .B0(n40), .B1(n894), .Y(n686) );
  CMPR42X1 U1617 ( .A(n797), .B(n702), .C(n759), .D(n740), .ICI(n563), .S(n556), .ICO(n554), .CO(n555) );
  OAI22XL U1618 ( .A0(n29), .A1(n949), .B0(n27), .B1(n948), .Y(n740) );
  OAI22XL U1619 ( .A0(n23), .A1(n968), .B0(n21), .B1(n967), .Y(n759) );
  OAI22XL U1620 ( .A0(n41), .A1(n911), .B0(n40), .B1(n910), .Y(n702) );
  CMPR42X1 U1621 ( .A(n693), .B(n459), .C(n456), .D(n460), .ICI(n457), .S(n442), .ICO(n440), .CO(n441) );
  OAI22XL U1622 ( .A0(n1073), .A1(n902), .B0(n40), .B1(n901), .Y(n693) );
  CMPR42X1 U1623 ( .A(n675), .B(n656), .C(n472), .D(n469), .ICI(n458), .S(n455), .ICO(n453), .CO(n454) );
  OAI22XL U1624 ( .A0(n53), .A1(n865), .B0(n51), .B1(n864), .Y(n656) );
  OAI22XL U1625 ( .A0(n47), .A1(n884), .B0(n46), .B1(n883), .Y(n675) );
  NAND2X1 U1626 ( .A(n619), .B(n827), .Y(n299) );
  CMPR42X1 U1627 ( .A(n636), .B(n709), .C(n690), .D(n652), .ICI(n418), .S(n411), .ICO(n409), .CO(n410) );
  OAI22XL U1628 ( .A0(n53), .A1(n861), .B0(n51), .B1(n860), .Y(n652) );
  OAI22XL U1629 ( .A0(n1073), .A1(n899), .B0(n40), .B1(n898), .Y(n690) );
  OAI22XL U1630 ( .A0(n1070), .A1(n842), .B0(n57), .B1(n841), .Y(n636) );
  OAI22XL U1631 ( .A0(n1078), .A1(n1011), .B0(n9), .B1(n1010), .Y(n802) );
  CMPR42X1 U1632 ( .A(n791), .B(n677), .C(n772), .D(n715), .ICI(n496), .S(n484), .ICO(n482), .CO(n483) );
  OAI22XL U1633 ( .A0(n35), .A1(n924), .B0(n33), .B1(n923), .Y(n715) );
  OAI22XL U1634 ( .A0(n17), .A1(n981), .B0(n16), .B1(n980), .Y(n772) );
  OAI22XL U1635 ( .A0(n47), .A1(n886), .B0(n46), .B1(n885), .Y(n677) );
  CMPR42X1 U1636 ( .A(n733), .B(n790), .C(n771), .D(n752), .ICI(n482), .S(n470), .ICO(n468), .CO(n469) );
  OAI22XL U1637 ( .A0(n24), .A1(n961), .B0(n22), .B1(n960), .Y(n752) );
  OAI22XL U1638 ( .A0(n17), .A1(n980), .B0(n16), .B1(n979), .Y(n771) );
  OAI22XL U1639 ( .A0(n12), .A1(n999), .B0(n9), .B1(n998), .Y(n790) );
  CMPR42X1 U1640 ( .A(n474), .B(n770), .C(n751), .D(n789), .ICI(n471), .S(n461), .ICO(n459), .CO(n460) );
  AO21X1 U1641 ( .A0(n12), .A1(n9), .B0(n998), .Y(n789) );
  OAI22XL U1642 ( .A0(n24), .A1(n960), .B0(n22), .B1(n959), .Y(n751) );
  OAI22XL U1643 ( .A0(n17), .A1(n979), .B0(n16), .B1(n978), .Y(n770) );
  CMPR42X1 U1644 ( .A(n762), .B(n800), .C(n781), .D(n585), .ICI(n586), .S(n583), .ICO(n581), .CO(n582) );
  OAI22XL U1645 ( .A0(n17), .A1(n990), .B0(n15), .B1(n989), .Y(n781) );
  CMPR42X1 U1646 ( .A(n735), .B(n716), .C(n513), .D(n514), .ICI(n511), .S(n495), .ICO(n493), .CO(n494) );
  OAI22XL U1647 ( .A0(n35), .A1(n925), .B0(n33), .B1(n924), .Y(n716) );
  OAI22XL U1648 ( .A0(n30), .A1(n944), .B0(n27), .B1(n943), .Y(n735) );
  CMPR42X1 U1649 ( .A(n638), .B(n732), .C(n713), .D(n694), .ICI(n468), .S(n458), .ICO(n456), .CO(n457) );
  OAI22XL U1650 ( .A0(n41), .A1(n903), .B0(n1083), .B1(n902), .Y(n694) );
  OAI22XL U1651 ( .A0(n36), .A1(n922), .B0(n34), .B1(n921), .Y(n713) );
  OAI22XL U1652 ( .A0(n30), .A1(n941), .B0(n27), .B1(n940), .Y(n732) );
  ADDFXL U1653 ( .A(n712), .B(n769), .CI(n1225), .CO(n446), .S(n447) );
  OAI22XL U1654 ( .A0(n36), .A1(n921), .B0(n34), .B1(n920), .Y(n712) );
  OAI22XL U1655 ( .A0(n17), .A1(n978), .B0(n16), .B1(n977), .Y(n769) );
  ADDFXL U1656 ( .A(n448), .B(n749), .CI(n654), .CO(n435), .S(n436) );
  OAI22XL U1657 ( .A0(n53), .A1(n863), .B0(n51), .B1(n862), .Y(n654) );
  OAI22XL U1658 ( .A0(n24), .A1(n958), .B0(n22), .B1(n957), .Y(n749) );
  ADDFXL U1659 ( .A(n670), .B(n727), .CI(n405), .CO(n402), .S(n403) );
  OAI22XL U1660 ( .A0(n47), .A1(n879), .B0(n46), .B1(n878), .Y(n670) );
  CLKINVX1 U1661 ( .A(n1185), .Y(n405) );
  OAI22XL U1662 ( .A0(n41), .A1(n1209), .B0(n40), .B1(n913), .Y(n623) );
  OAI22XL U1663 ( .A0(n29), .A1(n950), .B0(n27), .B1(n949), .Y(n741) );
  OAI22XL U1664 ( .A0(n54), .A1(n1091), .B0(n51), .B1(n871), .Y(n621) );
  ADDFXL U1665 ( .A(n1185), .B(n707), .CI(n650), .CO(n394), .S(n395) );
  OAI22XL U1666 ( .A0(n54), .A1(n859), .B0(n51), .B1(n858), .Y(n650) );
  OAI22XL U1667 ( .A0(n36), .A1(n916), .B0(n34), .B1(n915), .Y(n707) );
  ADDFXL U1668 ( .A(n764), .B(n625), .CI(n783), .CO(n595), .S(n596) );
  OAI22X1 U1669 ( .A0(n1070), .A1(n835), .B0(n58), .B1(n834), .Y(n360) );
  CMPR42X1 U1670 ( .A(n664), .B(n645), .C(n361), .D(n365), .ICI(n362), .S(n359), .ICO(n357), .CO(n358) );
  OAI22XL U1671 ( .A0(n54), .A1(n854), .B0(n51), .B1(n853), .Y(n645) );
  OAI22XL U1672 ( .A0(n47), .A1(n873), .B0(n46), .B1(n872), .Y(n664) );
  CLKINVX1 U1673 ( .A(n360), .Y(n361) );
  CMPR42X1 U1674 ( .A(n633), .B(n684), .C(n366), .D(n370), .ICI(n367), .S(n364), .ICO(n362), .CO(n363) );
  AO21X1 U1675 ( .A0(n1073), .A1(n40), .B0(n893), .Y(n684) );
  OAI22XL U1676 ( .A0(n1070), .A1(n836), .B0(n58), .B1(n835), .Y(n633) );
  CMPR42X1 U1677 ( .A(n360), .B(n632), .C(n644), .D(n663), .ICI(n357), .S(n356), .ICO(n354), .CO(n355) );
  OAI22XL U1678 ( .A0(n54), .A1(n853), .B0(n51), .B1(n852), .Y(n644) );
  OAI22XL U1679 ( .A0(n1070), .A1(n834), .B0(n58), .B1(n833), .Y(n632) );
  OAI22XL U1680 ( .A0(n47), .A1(n874), .B0(n46), .B1(n873), .Y(n665) );
  OAI22XL U1681 ( .A0(n54), .A1(n855), .B0(n51), .B1(n854), .Y(n646) );
  ADDFXL U1682 ( .A(n647), .B(n666), .CI(n373), .CO(n370), .S(n371) );
  OAI22XL U1683 ( .A0(n54), .A1(n856), .B0(n51), .B1(n855), .Y(n647) );
  OAI22XL U1684 ( .A0(n47), .A1(n875), .B0(n46), .B1(n874), .Y(n666) );
  CLKINVX1 U1685 ( .A(n372), .Y(n373) );
  OAI22XL U1686 ( .A0(n1070), .A1(n833), .B0(n58), .B1(n832), .Y(n352) );
  OAI22XL U1687 ( .A0(n54), .A1(n852), .B0(n51), .B1(n851), .Y(n643) );
  CLKINVX1 U1688 ( .A(n352), .Y(n353) );
  OAI22XL U1689 ( .A0(n1070), .A1(n832), .B0(n58), .B1(n831), .Y(n631) );
  XNOR2X1 U1690 ( .A(n1239), .B(n61), .Y(n1038) );
  OAI22XL U1691 ( .A0(n5), .A1(n1033), .B0(n1032), .B1(n3), .Y(n824) );
  OAI22XL U1692 ( .A0(n1078), .A1(n1014), .B0(n9), .B1(n1013), .Y(n805) );
  OAI22XL U1693 ( .A0(n29), .A1(n952), .B0(n27), .B1(n951), .Y(n743) );
  CLKINVX1 U1694 ( .A(n31), .Y(n1094) );
  XNOR2X1 U1695 ( .A(n1239), .B(b[6]), .Y(n1032) );
  XNOR2X1 U1696 ( .A(n1239), .B(b[5]), .Y(n1033) );
  XNOR2X1 U1697 ( .A(n1239), .B(b[7]), .Y(n1031) );
  XNOR2X1 U1698 ( .A(n1239), .B(b[8]), .Y(n1030) );
  XNOR2X1 U1699 ( .A(n1239), .B(b[17]), .Y(n1021) );
  XNOR2X1 U1700 ( .A(n1239), .B(b[11]), .Y(n1027) );
  XNOR2X1 U1701 ( .A(n1239), .B(b[12]), .Y(n1026) );
  XNOR2X1 U1702 ( .A(n1239), .B(n1044), .Y(n1023) );
  XNOR2X1 U1703 ( .A(n1239), .B(b[14]), .Y(n1024) );
  XNOR2X1 U1704 ( .A(n1239), .B(n1046), .Y(n1025) );
  XNOR2X1 U1705 ( .A(n1239), .B(b[16]), .Y(n1022) );
  XNOR2X1 U1706 ( .A(n1239), .B(n1041), .Y(n1020) );
  XNOR2X1 U1707 ( .A(a[1]), .B(n1050), .Y(n1029) );
  XNOR2X1 U1708 ( .A(n1239), .B(n1049), .Y(n1028) );
  XNOR2X1 U1709 ( .A(n1239), .B(b[4]), .Y(n1034) );
  XNOR2X1 U1710 ( .A(n1239), .B(b[3]), .Y(n1035) );
  XNOR2X1 U1711 ( .A(n1233), .B(n1058), .Y(n995) );
  XNOR2X1 U1712 ( .A(n1205), .B(b[3]), .Y(n1014) );
  XNOR2X1 U1713 ( .A(n1205), .B(b[6]), .Y(n1011) );
  XNOR2X1 U1714 ( .A(n1241), .B(n1058), .Y(n974) );
  XNOR2X1 U1715 ( .A(n1205), .B(b[5]), .Y(n1012) );
  XNOR2X1 U1716 ( .A(n1205), .B(b[4]), .Y(n1013) );
  XNOR2X1 U1717 ( .A(n1233), .B(b[3]), .Y(n993) );
  XNOR2X1 U1718 ( .A(n1205), .B(b[11]), .Y(n1006) );
  XNOR2X1 U1719 ( .A(n31), .B(b[6]), .Y(n927) );
  XNOR2X1 U1720 ( .A(n31), .B(b[7]), .Y(n926) );
  XNOR2X1 U1721 ( .A(n1205), .B(b[14]), .Y(n1003) );
  XNOR2X1 U1722 ( .A(n1205), .B(n1044), .Y(n1002) );
  XNOR2X1 U1723 ( .A(n1245), .B(b[4]), .Y(n950) );
  XNOR2X1 U1724 ( .A(n1245), .B(b[3]), .Y(n951) );
  XNOR2X1 U1725 ( .A(n43), .B(n1058), .Y(n890) );
  XNOR2X1 U1726 ( .A(n1210), .B(b[3]), .Y(n909) );
  XNOR2X1 U1727 ( .A(n1241), .B(n1049), .Y(n965) );
  XNOR2X1 U1728 ( .A(n1233), .B(b[8]), .Y(n988) );
  XNOR2X1 U1729 ( .A(n1241), .B(b[11]), .Y(n964) );
  XNOR2X1 U1730 ( .A(n1241), .B(b[6]), .Y(n969) );
  XNOR2X1 U1731 ( .A(n31), .B(b[2]), .Y(n931) );
  XNOR2X1 U1732 ( .A(n1205), .B(n1046), .Y(n1004) );
  XNOR2X1 U1733 ( .A(n1245), .B(b[8]), .Y(n946) );
  XNOR2X1 U1734 ( .A(n1245), .B(b[7]), .Y(n947) );
  XNOR2X1 U1735 ( .A(n1233), .B(b[11]), .Y(n985) );
  XNOR2X1 U1736 ( .A(n1241), .B(n1050), .Y(n966) );
  XNOR2X1 U1737 ( .A(n31), .B(b[5]), .Y(n928) );
  XNOR2X1 U1738 ( .A(n31), .B(b[4]), .Y(n929) );
  XNOR2X1 U1739 ( .A(n31), .B(b[3]), .Y(n930) );
  XNOR2X1 U1740 ( .A(n1233), .B(n1050), .Y(n987) );
  XNOR2X1 U1741 ( .A(n1233), .B(n1049), .Y(n986) );
  XNOR2X1 U1742 ( .A(n1205), .B(b[12]), .Y(n1005) );
  XNOR2X1 U1743 ( .A(n1210), .B(n1058), .Y(n911) );
  XNOR2X1 U1744 ( .A(n1210), .B(b[2]), .Y(n910) );
  XNOR2X1 U1745 ( .A(n1241), .B(b[8]), .Y(n967) );
  XNOR2X1 U1746 ( .A(n1241), .B(b[7]), .Y(n968) );
  XNOR2X1 U1747 ( .A(n1245), .B(b[5]), .Y(n949) );
  XNOR2X1 U1748 ( .A(n1245), .B(b[6]), .Y(n948) );
  XNOR2X1 U1749 ( .A(n31), .B(b[8]), .Y(n925) );
  XNOR2X1 U1750 ( .A(n1205), .B(b[16]), .Y(n1001) );
  XNOR2X1 U1751 ( .A(n1210), .B(b[6]), .Y(n906) );
  XNOR2X1 U1752 ( .A(n1241), .B(b[12]), .Y(n963) );
  XNOR2X1 U1753 ( .A(n1241), .B(n1046), .Y(n962) );
  XNOR2X1 U1754 ( .A(n43), .B(b[4]), .Y(n887) );
  XNOR2X1 U1755 ( .A(n1205), .B(b[17]), .Y(n1000) );
  XNOR2X1 U1756 ( .A(n43), .B(b[5]), .Y(n886) );
  XNOR2X1 U1757 ( .A(n1233), .B(n1044), .Y(n981) );
  XNOR2X1 U1758 ( .A(n31), .B(n1050), .Y(n924) );
  XNOR2X1 U1759 ( .A(n1216), .B(b[2]), .Y(n847) );
  XNOR2X1 U1760 ( .A(n1216), .B(n1058), .Y(n848) );
  XNOR2X1 U1761 ( .A(n1245), .B(b[12]), .Y(n942) );
  XNOR2X1 U1762 ( .A(n1245), .B(b[11]), .Y(n943) );
  XNOR2X1 U1763 ( .A(n1210), .B(b[7]), .Y(n905) );
  XNOR2X1 U1764 ( .A(n1183), .B(b[3]), .Y(n867) );
  XNOR2X1 U1765 ( .A(n1183), .B(n1058), .Y(n869) );
  XNOR2X1 U1766 ( .A(n1183), .B(b[2]), .Y(n868) );
  XNOR2X1 U1767 ( .A(n1233), .B(b[14]), .Y(n982) );
  XNOR2X1 U1768 ( .A(n1245), .B(n1049), .Y(n944) );
  XNOR2X1 U1769 ( .A(n1245), .B(n1050), .Y(n945) );
  XNOR2X1 U1770 ( .A(n1233), .B(b[12]), .Y(n984) );
  XNOR2X1 U1771 ( .A(n1233), .B(n1046), .Y(n983) );
  XNOR2X1 U1772 ( .A(n43), .B(b[3]), .Y(n888) );
  XNOR2X1 U1773 ( .A(n43), .B(b[2]), .Y(n889) );
  XNOR2X1 U1774 ( .A(n1210), .B(b[4]), .Y(n908) );
  XNOR2X1 U1775 ( .A(n1210), .B(b[5]), .Y(n907) );
  XNOR2X1 U1776 ( .A(n1216), .B(b[4]), .Y(n845) );
  XNOR2X1 U1777 ( .A(n1216), .B(b[5]), .Y(n844) );
  XNOR2X1 U1778 ( .A(n31), .B(n1049), .Y(n923) );
  XNOR2X1 U1779 ( .A(n43), .B(b[6]), .Y(n885) );
  XNOR2X1 U1780 ( .A(n1205), .B(n1041), .Y(n999) );
  XNOR2X1 U1781 ( .A(n1233), .B(b[16]), .Y(n980) );
  XNOR2X1 U1782 ( .A(n1241), .B(b[14]), .Y(n961) );
  XNOR2X1 U1783 ( .A(n1210), .B(b[8]), .Y(n904) );
  XNOR2X1 U1784 ( .A(n1183), .B(b[5]), .Y(n865) );
  XNOR2X1 U1785 ( .A(n1183), .B(b[4]), .Y(n866) );
  XNOR2X1 U1786 ( .A(n1233), .B(b[17]), .Y(n979) );
  XNOR2X1 U1787 ( .A(n1241), .B(b[16]), .Y(n959) );
  XNOR2X1 U1788 ( .A(n1241), .B(n1044), .Y(n960) );
  XNOR2X1 U1789 ( .A(n1216), .B(b[3]), .Y(n846) );
  XNOR2X1 U1790 ( .A(n1245), .B(n1046), .Y(n941) );
  XNOR2X1 U1791 ( .A(n31), .B(b[11]), .Y(n922) );
  XNOR2X1 U1792 ( .A(n1210), .B(n1050), .Y(n903) );
  XNOR2X1 U1793 ( .A(n1210), .B(n1049), .Y(n902) );
  XNOR2X1 U1794 ( .A(n1233), .B(n1041), .Y(n978) );
  XNOR2X1 U1795 ( .A(n31), .B(b[12]), .Y(n921) );
  XNOR2X1 U1796 ( .A(n31), .B(n1046), .Y(n920) );
  XNOR2X1 U1797 ( .A(n1241), .B(b[17]), .Y(n958) );
  XNOR2X1 U1798 ( .A(n1183), .B(b[7]), .Y(n863) );
  XNOR2X1 U1799 ( .A(n1183), .B(b[6]), .Y(n864) );
  XNOR2X1 U1800 ( .A(n1245), .B(b[14]), .Y(n940) );
  XNOR2X1 U1801 ( .A(n1245), .B(n1044), .Y(n939) );
  XNOR2X1 U1802 ( .A(n1216), .B(b[6]), .Y(n843) );
  XNOR2X1 U1803 ( .A(n1216), .B(b[7]), .Y(n842) );
  XNOR2X1 U1804 ( .A(n1216), .B(n1049), .Y(n839) );
  XNOR2X1 U1805 ( .A(n1216), .B(b[11]), .Y(n838) );
  XNOR2X1 U1806 ( .A(n1241), .B(b[2]), .Y(n973) );
  XNOR2X1 U1807 ( .A(n1233), .B(b[4]), .Y(n992) );
  XNOR2X1 U1808 ( .A(n13), .B(b[5]), .Y(n991) );
  XNOR2X1 U1809 ( .A(n1241), .B(b[3]), .Y(n972) );
  XNOR2X1 U1810 ( .A(n1205), .B(b[7]), .Y(n1010) );
  XNOR2X1 U1811 ( .A(n31), .B(n1058), .Y(n932) );
  XNOR2X1 U1812 ( .A(n1205), .B(b[2]), .Y(n1015) );
  XNOR2X1 U1813 ( .A(n1205), .B(n1058), .Y(n1016) );
  XNOR2X1 U1814 ( .A(n1245), .B(n1058), .Y(n953) );
  XNOR2X1 U1815 ( .A(n1245), .B(b[2]), .Y(n952) );
  XNOR2X1 U1816 ( .A(n1241), .B(b[5]), .Y(n970) );
  XNOR2X1 U1817 ( .A(n1241), .B(b[4]), .Y(n971) );
  XNOR2X1 U1818 ( .A(n1205), .B(b[8]), .Y(n1009) );
  XNOR2X1 U1819 ( .A(n1233), .B(b[7]), .Y(n989) );
  XNOR2X1 U1820 ( .A(n1233), .B(b[6]), .Y(n990) );
  XNOR2X1 U1821 ( .A(n1239), .B(n1040), .Y(n1019) );
  XNOR2X1 U1822 ( .A(n1205), .B(n1040), .Y(n998) );
  XNOR2X1 U1823 ( .A(n1233), .B(n1040), .Y(n977) );
  ADDHX1 U1824 ( .A(n628), .B(n808), .CO(n618), .S(n619) );
  OAI22XL U1825 ( .A0(n12), .A1(n1098), .B0(n9), .B1(n1018), .Y(n628) );
  XNOR2X1 U1826 ( .A(n1205), .B(n61), .Y(n1017) );
  XNOR2X1 U1827 ( .A(n1241), .B(n61), .Y(n975) );
  XNOR2X1 U1828 ( .A(n1216), .B(n61), .Y(n849) );
  ADDFX2 U1829 ( .A(n806), .B(n787), .CI(n615), .CO(n612), .S(n613) );
  OAI22XL U1830 ( .A0(n1078), .A1(n1015), .B0(n9), .B1(n1014), .Y(n806) );
  OAI22XL U1831 ( .A0(n17), .A1(n996), .B0(n15), .B1(n995), .Y(n787) );
  XNOR2X1 U1832 ( .A(n1233), .B(n61), .Y(n996) );
  ADDFX2 U1833 ( .A(n788), .B(n807), .CI(n826), .CO(n616), .S(n617) );
  OAI22XL U1834 ( .A0(n5), .A1(n1035), .B0(n1034), .B1(n3), .Y(n826) );
  NOR2BX1 U1835 ( .AN(n61), .B(n15), .Y(n788) );
  OAI22XL U1836 ( .A0(n1078), .A1(n1016), .B0(n9), .B1(n1015), .Y(n807) );
  OAI22XL U1837 ( .A0(n29), .A1(n954), .B0(n27), .B1(n953), .Y(n745) );
  XNOR2X1 U1838 ( .A(n1245), .B(n61), .Y(n954) );
  OAI22XL U1839 ( .A0(n41), .A1(n912), .B0(n40), .B1(n911), .Y(n703) );
  XNOR2X1 U1840 ( .A(n1210), .B(n61), .Y(n912) );
  XNOR2X1 U1841 ( .A(n1183), .B(n61), .Y(n870) );
  XNOR2X1 U1842 ( .A(n31), .B(n61), .Y(n933) );
  NOR2BX1 U1843 ( .AN(n61), .B(n46), .Y(n683) );
  OAI22XL U1844 ( .A0(n17), .A1(n987), .B0(n15), .B1(n986), .Y(n778) );
  CMPR42X1 U1845 ( .A(n641), .B(n679), .C(n755), .D(n812), .ICI(n525), .S(n515), .ICO(n513), .CO(n514) );
  OAI22XL U1846 ( .A0(n5), .A1(n1021), .B0(n1020), .B1(n3), .Y(n812) );
  NOR2BX1 U1847 ( .AN(n61), .B(n57), .Y(n641) );
  OAI22XL U1848 ( .A0(n24), .A1(n964), .B0(n22), .B1(n963), .Y(n755) );
  OAI22XL U1849 ( .A0(n5), .A1(n1029), .B0(n1028), .B1(n3), .Y(n820) );
  NAND2BX1 U1850 ( .AN(n61), .B(n1241), .Y(n976) );
  NAND2BX1 U1851 ( .AN(n61), .B(n1210), .Y(n913) );
  NAND2BX1 U1852 ( .AN(n61), .B(n1183), .Y(n871) );
  NAND2BX1 U1853 ( .AN(n61), .B(n43), .Y(n892) );
  NAND2BX1 U1854 ( .AN(n61), .B(n1245), .Y(n955) );
  NAND2BX1 U1855 ( .AN(n61), .B(n1205), .Y(n1018) );
  NAND2BX1 U1856 ( .AN(n61), .B(n31), .Y(n934) );
  CLKBUFX3 U1857 ( .A(n1237), .Y(n22) );
  CLKBUFX3 U1858 ( .A(n1084), .Y(n34) );
  CLKBUFX3 U1859 ( .A(n1071), .Y(n54) );
  OAI22XL U1860 ( .A0(n23), .A1(n974), .B0(n21), .B1(n973), .Y(n765) );
  NOR2BX1 U1861 ( .AN(n61), .B(n51), .Y(n662) );
  OAI22XL U1862 ( .A0(n23), .A1(n966), .B0(n21), .B1(n965), .Y(n757) );
  OAI22XL U1863 ( .A0(n17), .A1(n989), .B0(n15), .B1(n988), .Y(n780) );
  CLKINVX1 U1864 ( .A(n1183), .Y(n1091) );
  CLKINVX1 U1865 ( .A(n43), .Y(n1092) );
  XNOR2X1 U1866 ( .A(n43), .B(b[7]), .Y(n884) );
  XNOR2X1 U1867 ( .A(n1210), .B(b[11]), .Y(n901) );
  XNOR2X1 U1868 ( .A(n43), .B(b[8]), .Y(n883) );
  XNOR2X1 U1869 ( .A(n43), .B(n1050), .Y(n882) );
  XNOR2X1 U1870 ( .A(n1210), .B(b[12]), .Y(n900) );
  XNOR2X1 U1871 ( .A(n1241), .B(n1041), .Y(n957) );
  XNOR2X1 U1872 ( .A(n1183), .B(b[8]), .Y(n862) );
  XNOR2X1 U1873 ( .A(n1210), .B(n1046), .Y(n899) );
  XNOR2X1 U1874 ( .A(n1183), .B(n1050), .Y(n861) );
  XNOR2X1 U1875 ( .A(n1245), .B(b[17]), .Y(n937) );
  XNOR2X1 U1876 ( .A(n1245), .B(b[16]), .Y(n938) );
  XNOR2X1 U1877 ( .A(n43), .B(n1049), .Y(n881) );
  XNOR2X1 U1878 ( .A(n43), .B(b[11]), .Y(n880) );
  XNOR2X1 U1879 ( .A(n31), .B(n1044), .Y(n918) );
  XNOR2X1 U1880 ( .A(n31), .B(b[14]), .Y(n919) );
  XNOR2X1 U1881 ( .A(n1216), .B(n1050), .Y(n840) );
  XNOR2X1 U1882 ( .A(n1216), .B(b[8]), .Y(n841) );
  XNOR2X1 U1883 ( .A(n1183), .B(b[12]), .Y(n858) );
  XNOR2X1 U1884 ( .A(n1245), .B(n1041), .Y(n936) );
  XNOR2X1 U1885 ( .A(n43), .B(b[12]), .Y(n879) );
  XNOR2X1 U1886 ( .A(n1216), .B(n1046), .Y(n836) );
  XNOR2X1 U1887 ( .A(n1216), .B(b[12]), .Y(n837) );
  XNOR2X1 U1888 ( .A(n31), .B(b[17]), .Y(n916) );
  XNOR2X1 U1889 ( .A(n31), .B(b[16]), .Y(n917) );
  XNOR2X1 U1890 ( .A(n1183), .B(b[11]), .Y(n859) );
  XNOR2X1 U1891 ( .A(n1183), .B(n1049), .Y(n860) );
  XNOR2X1 U1892 ( .A(n1210), .B(b[14]), .Y(n898) );
  XNOR2X1 U1893 ( .A(n31), .B(n1041), .Y(n915) );
  XNOR2X1 U1894 ( .A(n1210), .B(b[16]), .Y(n896) );
  XNOR2X1 U1895 ( .A(n1210), .B(n1044), .Y(n897) );
  XNOR2X1 U1896 ( .A(n43), .B(b[14]), .Y(n877) );
  XNOR2X1 U1897 ( .A(n43), .B(n1046), .Y(n878) );
  XNOR2X1 U1898 ( .A(n43), .B(b[17]), .Y(n874) );
  XNOR2X1 U1899 ( .A(n1183), .B(n1044), .Y(n855) );
  XNOR2X1 U1900 ( .A(n1183), .B(b[14]), .Y(n856) );
  XNOR2X1 U1901 ( .A(n1210), .B(b[17]), .Y(n895) );
  XNOR2X1 U1902 ( .A(n43), .B(n1044), .Y(n876) );
  XNOR2X1 U1903 ( .A(n43), .B(b[16]), .Y(n875) );
  XNOR2X1 U1904 ( .A(n1183), .B(n1046), .Y(n857) );
  XNOR2X1 U1905 ( .A(n1210), .B(n1041), .Y(n894) );
  XNOR2X1 U1906 ( .A(n43), .B(n1041), .Y(n873) );
  XNOR2X1 U1907 ( .A(n1183), .B(b[16]), .Y(n854) );
  XNOR2X1 U1908 ( .A(n1216), .B(b[14]), .Y(n835) );
  XNOR2X1 U1909 ( .A(n1216), .B(n1044), .Y(n834) );
  XNOR2X1 U1910 ( .A(n1183), .B(b[17]), .Y(n853) );
  XNOR2X1 U1911 ( .A(n1241), .B(n1040), .Y(n956) );
  XNOR2X1 U1912 ( .A(n1245), .B(n1040), .Y(n935) );
  XNOR2X1 U1913 ( .A(n31), .B(n1040), .Y(n914) );
  XNOR2X1 U1914 ( .A(n1210), .B(n1040), .Y(n893) );
  XNOR2X1 U1915 ( .A(n43), .B(n1040), .Y(n872) );
  CLKINVX1 U1916 ( .A(n1205), .Y(n1098) );
  XNOR2X1 U1917 ( .A(n1216), .B(b[17]), .Y(n832) );
  XNOR2X1 U1918 ( .A(n1216), .B(b[16]), .Y(n833) );
  XNOR2X1 U1919 ( .A(n1183), .B(n1041), .Y(n852) );
  XNOR2X1 U1920 ( .A(n1216), .B(n1041), .Y(n831) );
  XNOR2X1 U1921 ( .A(n1183), .B(n1040), .Y(n851) );
  XNOR2X1 U1922 ( .A(n1216), .B(n1040), .Y(n830) );
  XOR2X1 U1923 ( .A(a[13]), .B(a[12]), .Y(n1063) );
  XOR2X1 U1924 ( .A(a[7]), .B(a[6]), .Y(n1066) );
  XOR2X1 U1925 ( .A(a[19]), .B(a[18]), .Y(n1060) );
  XOR2X1 U1926 ( .A(a[17]), .B(a[16]), .Y(n1061) );
  XOR2X1 U1927 ( .A(a[9]), .B(a[8]), .Y(n1065) );
  XOR2X1 U1928 ( .A(a[11]), .B(a[10]), .Y(n1064) );
  XOR2X1 U1929 ( .A(a[3]), .B(a[2]), .Y(n1068) );
  NAND2X1 U1930 ( .A(n1069), .B(n1089), .Y(n1079) );
  XOR2X1 U1931 ( .A(a[0]), .B(a[1]), .Y(n1069) );
endmodule


module CONV_DW01_add_8 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n55, n57, n58, n59, n60, n61,
         n62, n63, n64, n66, n68, n69, n70, n72, n73, n74, n75, n76, n77, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n116, n118, n120, n121,
         n122, n123, n125, n126, n128, n129, n130, n131, n132, n134, n136,
         n137, n138, n141, n143, n144, n145, n146, n147, n149, n151, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n172, n174, n175, n176, n179,
         n181, n182, n183, n184, n185, n187, n189, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n220, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n238, n240, n241, n242,
         n243, n244, n246, n248, n249, n250, n251, n252, n254, n256, n257,
         n258, n259, n260, n261, n263, n264, n269, n270, n271, n272, n273,
         n274, n277, n281, n283, n288, n289, n296, n298, n300, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456;

  XNOR2X2 U345 ( .A(n58), .B(n4), .Y(SUM[36]) );
  XNOR2X2 U346 ( .A(n51), .B(n3), .Y(SUM[37]) );
  NAND2X1 U347 ( .A(B[8]), .B(A[8]), .Y(n229) );
  NOR2X4 U348 ( .A(n440), .B(n445), .Y(n76) );
  NAND2X1 U349 ( .A(n85), .B(n93), .Y(n83) );
  NAND2X1 U350 ( .A(n447), .B(n64), .Y(n62) );
  AOI21X1 U351 ( .A0(n430), .A1(n73), .B0(n66), .Y(n64) );
  CLKINVX1 U352 ( .A(n68), .Y(n66) );
  NOR2X1 U353 ( .A(B[20]), .B(A[20]), .Y(n155) );
  OR2X1 U354 ( .A(B[16]), .B(A[16]), .Y(n435) );
  CLKINVX1 U355 ( .A(n194), .Y(n192) );
  OR2X1 U356 ( .A(B[15]), .B(A[15]), .Y(n433) );
  CLKINVX1 U357 ( .A(n136), .Y(n134) );
  OR2X1 U358 ( .A(B[35]), .B(A[35]), .Y(n430) );
  OR2X1 U359 ( .A(n81), .B(n52), .Y(n442) );
  CLKINVX1 U360 ( .A(n174), .Y(n172) );
  OR2X1 U361 ( .A(B[26]), .B(A[26]), .Y(n432) );
  OR2X4 U362 ( .A(n81), .B(n59), .Y(n443) );
  OR2X1 U363 ( .A(B[36]), .B(A[36]), .Y(n431) );
  OR2X1 U364 ( .A(B[17]), .B(A[17]), .Y(n429) );
  OR2X1 U365 ( .A(B[22]), .B(A[22]), .Y(n444) );
  OR2X1 U366 ( .A(B[21]), .B(A[21]), .Y(n428) );
  OR2X1 U367 ( .A(B[2]), .B(A[2]), .Y(n438) );
  OR2X1 U368 ( .A(B[4]), .B(A[4]), .Y(n437) );
  CLKINVX1 U369 ( .A(n234), .Y(n232) );
  OR2X1 U370 ( .A(B[23]), .B(A[23]), .Y(n434) );
  CLKINVX1 U371 ( .A(n216), .Y(n214) );
  NAND2X1 U372 ( .A(B[12]), .B(A[12]), .Y(n203) );
  NOR2X1 U373 ( .A(B[12]), .B(A[12]), .Y(n202) );
  NAND2X1 U374 ( .A(B[27]), .B(A[27]), .Y(n110) );
  XOR2X1 U375 ( .A(n76), .B(n6), .Y(SUM[34]) );
  XOR2X1 U376 ( .A(n81), .B(n7), .Y(SUM[33]) );
  XOR2X1 U377 ( .A(n46), .B(n2), .Y(SUM[38]) );
  NAND2XL U378 ( .A(n72), .B(n75), .Y(n6) );
  OAI21X4 U379 ( .A0(n76), .A1(n70), .B0(n75), .Y(n69) );
  NAND2X1 U380 ( .A(B[34]), .B(A[34]), .Y(n75) );
  OR2X1 U381 ( .A(B[9]), .B(A[9]), .Y(n436) );
  OR2X1 U382 ( .A(B[6]), .B(A[6]), .Y(n439) );
  NAND2X1 U383 ( .A(B[21]), .B(A[21]), .Y(n151) );
  NAND2X1 U384 ( .A(B[33]), .B(A[33]), .Y(n80) );
  CLKINVX1 U385 ( .A(n80), .Y(n445) );
  NAND2X1 U386 ( .A(B[22]), .B(A[22]), .Y(n143) );
  NOR2X1 U387 ( .A(B[33]), .B(A[33]), .Y(n79) );
  CLKINVX1 U388 ( .A(n193), .Y(n191) );
  NAND2X1 U389 ( .A(B[16]), .B(A[16]), .Y(n181) );
  CLKINVX1 U390 ( .A(n215), .Y(n213) );
  CLKINVX1 U391 ( .A(n233), .Y(n231) );
  CLKINVX1 U392 ( .A(n210), .Y(n208) );
  OAI21X1 U393 ( .A0(n53), .A1(n49), .B0(n50), .Y(n48) );
  AOI21X2 U394 ( .A0(n223), .A1(n436), .B0(n220), .Y(n218) );
  NOR2X1 U395 ( .A(n95), .B(n100), .Y(n93) );
  NOR2X1 U396 ( .A(B[30]), .B(A[30]), .Y(n95) );
  INVXL U397 ( .A(n205), .Y(n204) );
  AOI21X4 U398 ( .A0(n197), .A1(n205), .B0(n198), .Y(n196) );
  OAI21X2 U399 ( .A0(n206), .A1(n218), .B0(n207), .Y(n205) );
  CLKINVX2 U400 ( .A(n82), .Y(n81) );
  AOI21X2 U401 ( .A0(n102), .A1(n93), .B0(n94), .Y(n92) );
  XOR2XL U402 ( .A(n92), .B(n9), .Y(SUM[31]) );
  AND2X1 U403 ( .A(n82), .B(n77), .Y(n440) );
  INVXL U404 ( .A(n79), .Y(n77) );
  XNOR2X4 U405 ( .A(n69), .B(n5), .Y(SUM[35]) );
  AND2X1 U406 ( .A(n82), .B(n47), .Y(n441) );
  NOR2X4 U407 ( .A(n441), .B(n48), .Y(n46) );
  NAND2X6 U408 ( .A(n455), .B(n84), .Y(n82) );
  OAI21X2 U409 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NAND2X1 U410 ( .A(n61), .B(n431), .Y(n52) );
  OAI21X1 U411 ( .A0(n95), .A1(n101), .B0(n96), .Y(n94) );
  AOI21X2 U412 ( .A0(n62), .A1(n431), .B0(n55), .Y(n53) );
  NAND2X1 U413 ( .A(B[26]), .B(A[26]), .Y(n118) );
  NAND2X1 U414 ( .A(B[15]), .B(A[15]), .Y(n189) );
  NAND2X4 U415 ( .A(n442), .B(n53), .Y(n51) );
  NAND2X1 U416 ( .A(n443), .B(n60), .Y(n58) );
  NAND2X1 U417 ( .A(n77), .B(n80), .Y(n7) );
  INVXL U418 ( .A(n62), .Y(n60) );
  INVXL U419 ( .A(n61), .Y(n59) );
  NOR2X1 U420 ( .A(n448), .B(n165), .Y(n163) );
  NAND2XL U421 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2X2 U422 ( .A(n430), .B(n72), .Y(n63) );
  INVXL U423 ( .A(n163), .Y(n162) );
  OAI21X1 U424 ( .A0(n170), .A1(n166), .B0(n167), .Y(n165) );
  OAI21X1 U425 ( .A0(n199), .A1(n203), .B0(n200), .Y(n198) );
  NAND2X2 U426 ( .A(n445), .B(n446), .Y(n447) );
  INVX3 U427 ( .A(n63), .Y(n446) );
  INVX3 U428 ( .A(n449), .Y(n125) );
  OAI21X2 U429 ( .A0(n224), .A1(n236), .B0(n225), .Y(n223) );
  OAI21X2 U430 ( .A0(n244), .A1(n242), .B0(n243), .Y(n241) );
  OAI21X2 U431 ( .A0(n163), .A1(n146), .B0(n147), .Y(n145) );
  OAI21X2 U432 ( .A0(n196), .A1(n184), .B0(n185), .Y(n183) );
  OA21X4 U433 ( .A0(n132), .A1(n128), .B0(n129), .Y(n450) );
  NOR2X1 U434 ( .A(n87), .B(n90), .Y(n85) );
  AND2X2 U435 ( .A(n183), .B(n164), .Y(n448) );
  NOR2X1 U436 ( .A(B[13]), .B(A[13]), .Y(n199) );
  NOR2X1 U437 ( .A(B[28]), .B(A[28]), .Y(n106) );
  OAI21X1 U438 ( .A0(n92), .A1(n90), .B0(n91), .Y(n89) );
  NOR2X1 U439 ( .A(B[8]), .B(A[8]), .Y(n228) );
  NOR2X1 U440 ( .A(B[11]), .B(A[11]), .Y(n210) );
  NOR2X1 U441 ( .A(B[18]), .B(A[18]), .Y(n166) );
  NOR2X1 U442 ( .A(n169), .B(n166), .Y(n164) );
  NOR2X1 U443 ( .A(n79), .B(n63), .Y(n61) );
  AOI21X1 U444 ( .A0(n226), .A1(n232), .B0(n227), .Y(n225) );
  NAND2X1 U445 ( .A(n432), .B(n120), .Y(n113) );
  AOI21X1 U446 ( .A0(n85), .A1(n94), .B0(n86), .Y(n84) );
  OAI21X1 U447 ( .A0(n250), .A1(n252), .B0(n251), .Y(n249) );
  NOR2X2 U448 ( .A(n160), .B(n155), .Y(n153) );
  OAI21X1 U449 ( .A0(n258), .A1(n261), .B0(n259), .Y(n257) );
  INVX1 U450 ( .A(n44), .Y(n263) );
  NAND2X1 U451 ( .A(B[20]), .B(A[20]), .Y(n156) );
  NAND2X1 U452 ( .A(B[5]), .B(A[5]), .Y(n243) );
  NOR2X1 U453 ( .A(B[27]), .B(A[27]), .Y(n109) );
  OAI21XL U454 ( .A0(n111), .A1(n109), .B0(n110), .Y(n108) );
  NOR2X1 U455 ( .A(B[34]), .B(A[34]), .Y(n74) );
  NOR2X1 U456 ( .A(B[25]), .B(A[25]), .Y(n122) );
  OAI2BB1X4 U457 ( .A0N(n126), .A1N(n145), .B0(n450), .Y(n449) );
  INVXL U458 ( .A(n72), .Y(n70) );
  INVXL U459 ( .A(n444), .Y(n138) );
  INVXL U460 ( .A(n435), .Y(n176) );
  OAI21X2 U461 ( .A0(n155), .A1(n161), .B0(n156), .Y(n154) );
  OAI21X4 U462 ( .A0(n125), .A1(n113), .B0(n114), .Y(n112) );
  CLKINVX3 U463 ( .A(n123), .Y(n121) );
  INVXL U464 ( .A(n101), .Y(n99) );
  INVXL U465 ( .A(n95), .Y(n271) );
  INVXL U466 ( .A(n160), .Y(n158) );
  INVXL U467 ( .A(n161), .Y(n159) );
  INVXL U468 ( .A(n155), .Y(n281) );
  INVXL U469 ( .A(n87), .Y(n269) );
  NAND2XL U470 ( .A(n270), .B(n91), .Y(n9) );
  INVXL U471 ( .A(n90), .Y(n270) );
  XNOR2XL U472 ( .A(n102), .B(n11), .Y(SUM[29]) );
  NAND2XL U473 ( .A(n272), .B(n101), .Y(n11) );
  INVXL U474 ( .A(n100), .Y(n272) );
  NAND2XL U475 ( .A(n274), .B(n110), .Y(n13) );
  INVXL U476 ( .A(n109), .Y(n274) );
  XNOR2X1 U477 ( .A(n451), .B(n10), .Y(SUM[30]) );
  AO21XL U478 ( .A0(n102), .A1(n272), .B0(n99), .Y(n451) );
  NOR2X1 U479 ( .A(B[24]), .B(A[24]), .Y(n128) );
  NAND2XL U480 ( .A(B[30]), .B(A[30]), .Y(n96) );
  NAND2XL U481 ( .A(B[24]), .B(A[24]), .Y(n129) );
  NAND2XL U482 ( .A(B[28]), .B(A[28]), .Y(n107) );
  NAND2XL U483 ( .A(B[32]), .B(A[32]), .Y(n88) );
  NAND2XL U484 ( .A(B[13]), .B(A[13]), .Y(n200) );
  NAND2XL U485 ( .A(n434), .B(n136), .Y(n17) );
  XNOR2X1 U486 ( .A(n452), .B(n19), .Y(SUM[21]) );
  AO21XL U487 ( .A0(n162), .A1(n153), .B0(n154), .Y(n452) );
  NAND2XL U488 ( .A(n281), .B(n156), .Y(n20) );
  XNOR2X1 U489 ( .A(n453), .B(n14), .Y(SUM[26]) );
  AO21XL U490 ( .A0(n449), .A1(n120), .B0(n121), .Y(n453) );
  NAND2XL U491 ( .A(n120), .B(n123), .Y(n15) );
  NAND2XL U492 ( .A(n444), .B(n143), .Y(n18) );
  NAND2XL U493 ( .A(n158), .B(n161), .Y(n21) );
  NOR2X1 U494 ( .A(B[37]), .B(A[37]), .Y(n49) );
  NAND2XL U495 ( .A(B[35]), .B(A[35]), .Y(n68) );
  NAND2XL U496 ( .A(B[37]), .B(A[37]), .Y(n50) );
  NAND2XL U497 ( .A(B[38]), .B(A[38]), .Y(n45) );
  NAND2XL U498 ( .A(B[39]), .B(A[39]), .Y(n42) );
  NAND2XL U499 ( .A(n435), .B(n181), .Y(n24) );
  NAND2XL U500 ( .A(n429), .B(n174), .Y(n23) );
  NAND2XL U501 ( .A(n283), .B(n167), .Y(n22) );
  NAND2XL U502 ( .A(n288), .B(n200), .Y(n27) );
  NAND2XL U503 ( .A(n213), .B(n216), .Y(n30) );
  NAND2XL U504 ( .A(n208), .B(n211), .Y(n29) );
  AOI21XL U505 ( .A0(n217), .A1(n213), .B0(n214), .Y(n212) );
  XOR2XL U506 ( .A(n204), .B(n28), .Y(SUM[12]) );
  NAND2XL U507 ( .A(n289), .B(n203), .Y(n28) );
  INVXL U508 ( .A(n202), .Y(n289) );
  NAND2XL U509 ( .A(n191), .B(n194), .Y(n26) );
  XNOR2X1 U510 ( .A(n454), .B(n25), .Y(SUM[15]) );
  AO21XL U511 ( .A0(n195), .A1(n191), .B0(n192), .Y(n454) );
  NAND2XL U512 ( .A(n226), .B(n229), .Y(n32) );
  AOI21XL U513 ( .A0(n235), .A1(n231), .B0(n232), .Y(n230) );
  XNOR2XL U514 ( .A(n223), .B(n31), .Y(SUM[9]) );
  NAND2XL U515 ( .A(n436), .B(n222), .Y(n31) );
  XNOR2XL U516 ( .A(n34), .B(n241), .Y(SUM[6]) );
  NAND2XL U517 ( .A(n439), .B(n240), .Y(n34) );
  NAND2XL U518 ( .A(n231), .B(n234), .Y(n33) );
  XOR2XL U519 ( .A(n244), .B(n35), .Y(SUM[5]) );
  NAND2XL U520 ( .A(n296), .B(n243), .Y(n35) );
  INVXL U521 ( .A(n242), .Y(n296) );
  NAND2BXL U522 ( .AN(n260), .B(n261), .Y(n40) );
  XOR2XL U523 ( .A(n39), .B(n261), .Y(SUM[1]) );
  NAND2XL U524 ( .A(n300), .B(n259), .Y(n39) );
  INVXL U525 ( .A(n258), .Y(n300) );
  XNOR2XL U526 ( .A(n38), .B(n257), .Y(SUM[2]) );
  NAND2XL U527 ( .A(n438), .B(n256), .Y(n38) );
  XOR2XL U528 ( .A(n37), .B(n252), .Y(SUM[3]) );
  NAND2XL U529 ( .A(n298), .B(n251), .Y(n37) );
  INVXL U530 ( .A(n250), .Y(n298) );
  XNOR2XL U531 ( .A(n36), .B(n249), .Y(SUM[4]) );
  NAND2XL U532 ( .A(n437), .B(n248), .Y(n36) );
  NOR2XL U533 ( .A(B[0]), .B(A[0]), .Y(n260) );
  OR2X2 U534 ( .A(n103), .B(n83), .Y(n455) );
  AOI21X2 U535 ( .A0(n112), .A1(n104), .B0(n105), .Y(n103) );
  NAND2X1 U536 ( .A(n429), .B(n435), .Y(n169) );
  NAND2X1 U537 ( .A(n434), .B(n444), .Y(n131) );
  CLKINVX1 U538 ( .A(n103), .Y(n102) );
  CLKINVX1 U539 ( .A(n112), .Y(n111) );
  CLKINVX1 U540 ( .A(n183), .Y(n182) );
  CLKINVX1 U541 ( .A(n145), .Y(n144) );
  CLKINVX1 U542 ( .A(n196), .Y(n195) );
  CLKINVX1 U543 ( .A(n236), .Y(n235) );
  CLKINVX1 U544 ( .A(n218), .Y(n217) );
  NOR2X1 U545 ( .A(n199), .B(n202), .Y(n197) );
  NOR2X1 U546 ( .A(n128), .B(n131), .Y(n126) );
  NOR2X1 U547 ( .A(n106), .B(n109), .Y(n104) );
  OAI21XL U548 ( .A0(n106), .A1(n110), .B0(n107), .Y(n105) );
  AOI21X1 U549 ( .A0(n433), .A1(n192), .B0(n187), .Y(n185) );
  NAND2X1 U550 ( .A(n433), .B(n191), .Y(n184) );
  CLKINVX1 U551 ( .A(n189), .Y(n187) );
  AOI21X1 U552 ( .A0(n432), .A1(n121), .B0(n116), .Y(n114) );
  NAND2X1 U553 ( .A(n208), .B(n213), .Y(n206) );
  AOI21X1 U554 ( .A0(n208), .A1(n214), .B0(n209), .Y(n207) );
  NAND2X1 U555 ( .A(n153), .B(n428), .Y(n146) );
  AOI21X1 U556 ( .A0(n428), .A1(n154), .B0(n149), .Y(n147) );
  AOI21X1 U557 ( .A0(n241), .A1(n439), .B0(n238), .Y(n236) );
  CLKINVX1 U558 ( .A(n240), .Y(n238) );
  CLKINVX1 U559 ( .A(n222), .Y(n220) );
  AOI21X1 U560 ( .A0(n437), .A1(n249), .B0(n246), .Y(n244) );
  CLKINVX1 U561 ( .A(n248), .Y(n246) );
  NOR2X1 U562 ( .A(n52), .B(n49), .Y(n47) );
  AOI21X1 U563 ( .A0(n257), .A1(n438), .B0(n254), .Y(n252) );
  CLKINVX1 U564 ( .A(n256), .Y(n254) );
  AOI21X1 U565 ( .A0(n429), .A1(n179), .B0(n172), .Y(n170) );
  AOI21X1 U566 ( .A0(n434), .A1(n141), .B0(n134), .Y(n132) );
  CLKINVX1 U567 ( .A(n57), .Y(n55) );
  NAND2X1 U568 ( .A(n226), .B(n231), .Y(n224) );
  CLKINVX1 U569 ( .A(n229), .Y(n227) );
  OAI21XL U570 ( .A0(n87), .A1(n91), .B0(n88), .Y(n86) );
  CLKINVX1 U571 ( .A(n74), .Y(n72) );
  CLKINVX1 U572 ( .A(n228), .Y(n226) );
  CLKINVX1 U573 ( .A(n122), .Y(n120) );
  CLKINVX1 U574 ( .A(n75), .Y(n73) );
  CLKINVX1 U575 ( .A(n181), .Y(n179) );
  CLKINVX1 U576 ( .A(n143), .Y(n141) );
  CLKINVX1 U577 ( .A(n151), .Y(n149) );
  CLKINVX1 U578 ( .A(n49), .Y(n264) );
  CLKINVX1 U579 ( .A(n118), .Y(n116) );
  CLKINVX1 U580 ( .A(n211), .Y(n209) );
  CLKINVX1 U581 ( .A(n106), .Y(n273) );
  CLKINVX1 U582 ( .A(n128), .Y(n277) );
  CLKINVX1 U583 ( .A(n199), .Y(n288) );
  CLKINVX1 U584 ( .A(n166), .Y(n283) );
  NOR2X1 U585 ( .A(B[29]), .B(A[29]), .Y(n100) );
  NOR2X1 U586 ( .A(B[19]), .B(A[19]), .Y(n160) );
  NOR2X1 U587 ( .A(B[31]), .B(A[31]), .Y(n90) );
  NOR2X2 U588 ( .A(B[32]), .B(A[32]), .Y(n87) );
  NOR2X1 U589 ( .A(B[7]), .B(A[7]), .Y(n233) );
  NOR2X1 U590 ( .A(B[10]), .B(A[10]), .Y(n215) );
  NOR2X1 U591 ( .A(B[14]), .B(A[14]), .Y(n193) );
  NOR2X1 U592 ( .A(B[38]), .B(A[38]), .Y(n44) );
  NOR2X1 U593 ( .A(B[5]), .B(A[5]), .Y(n242) );
  NOR2X1 U594 ( .A(B[1]), .B(A[1]), .Y(n258) );
  NOR2X1 U595 ( .A(B[3]), .B(A[3]), .Y(n250) );
  NAND2X1 U596 ( .A(n431), .B(n57), .Y(n4) );
  NAND2X1 U597 ( .A(B[29]), .B(A[29]), .Y(n101) );
  NAND2X1 U598 ( .A(B[31]), .B(A[31]), .Y(n91) );
  NAND2X1 U599 ( .A(B[19]), .B(A[19]), .Y(n161) );
  XNOR2X1 U600 ( .A(n89), .B(n8), .Y(SUM[32]) );
  NAND2X1 U601 ( .A(n269), .B(n88), .Y(n8) );
  NAND2X1 U602 ( .A(n430), .B(n68), .Y(n5) );
  NAND2X1 U603 ( .A(B[2]), .B(A[2]), .Y(n256) );
  NAND2X1 U604 ( .A(B[9]), .B(A[9]), .Y(n222) );
  NAND2X1 U605 ( .A(B[17]), .B(A[17]), .Y(n174) );
  NAND2X1 U606 ( .A(B[23]), .B(A[23]), .Y(n136) );
  NAND2X1 U607 ( .A(B[25]), .B(A[25]), .Y(n123) );
  NAND2X1 U608 ( .A(B[36]), .B(A[36]), .Y(n57) );
  NAND2X1 U609 ( .A(B[18]), .B(A[18]), .Y(n167) );
  NAND2X1 U610 ( .A(n432), .B(n118), .Y(n14) );
  XNOR2X1 U611 ( .A(n108), .B(n12), .Y(SUM[28]) );
  NAND2X1 U612 ( .A(n273), .B(n107), .Y(n12) );
  NAND2X1 U613 ( .A(n271), .B(n96), .Y(n10) );
  NAND2X1 U614 ( .A(n264), .B(n50), .Y(n3) );
  NAND2X1 U615 ( .A(n263), .B(n45), .Y(n2) );
  XNOR2X1 U616 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NAND2X1 U617 ( .A(n456), .B(n42), .Y(n1) );
  NAND2X1 U618 ( .A(B[4]), .B(A[4]), .Y(n248) );
  NAND2X1 U619 ( .A(B[6]), .B(A[6]), .Y(n240) );
  NAND2X1 U620 ( .A(B[7]), .B(A[7]), .Y(n234) );
  NAND2X1 U621 ( .A(B[10]), .B(A[10]), .Y(n216) );
  NAND2X1 U622 ( .A(B[14]), .B(A[14]), .Y(n194) );
  NAND2X1 U623 ( .A(B[1]), .B(A[1]), .Y(n259) );
  NAND2X1 U624 ( .A(B[3]), .B(A[3]), .Y(n251) );
  XOR2X1 U625 ( .A(n111), .B(n13), .Y(SUM[27]) );
  OR2X1 U626 ( .A(B[39]), .B(A[39]), .Y(n456) );
  XNOR2X1 U627 ( .A(n175), .B(n23), .Y(SUM[17]) );
  OAI21XL U628 ( .A0(n182), .A1(n176), .B0(n181), .Y(n175) );
  XNOR2X1 U629 ( .A(n137), .B(n17), .Y(SUM[23]) );
  OAI21XL U630 ( .A0(n144), .A1(n138), .B0(n143), .Y(n137) );
  XNOR2X1 U631 ( .A(n449), .B(n15), .Y(SUM[25]) );
  NAND2X1 U632 ( .A(n433), .B(n189), .Y(n25) );
  NAND2X1 U633 ( .A(B[0]), .B(A[0]), .Y(n261) );
  CLKINVX1 U634 ( .A(n40), .Y(SUM[0]) );
  XNOR2X1 U635 ( .A(n33), .B(n235), .Y(SUM[7]) );
  XOR2X1 U636 ( .A(n230), .B(n32), .Y(SUM[8]) );
  XNOR2X1 U637 ( .A(n217), .B(n30), .Y(SUM[10]) );
  XOR2X1 U638 ( .A(n212), .B(n29), .Y(SUM[11]) );
  XNOR2X1 U639 ( .A(n201), .B(n27), .Y(SUM[13]) );
  OAI21XL U640 ( .A0(n204), .A1(n202), .B0(n203), .Y(n201) );
  XNOR2X1 U641 ( .A(n195), .B(n26), .Y(SUM[14]) );
  XOR2X1 U642 ( .A(n182), .B(n24), .Y(SUM[16]) );
  XNOR2X1 U643 ( .A(n168), .B(n22), .Y(SUM[18]) );
  OAI21XL U644 ( .A0(n182), .A1(n169), .B0(n170), .Y(n168) );
  XNOR2X1 U645 ( .A(n162), .B(n21), .Y(SUM[19]) );
  XOR2X1 U646 ( .A(n157), .B(n20), .Y(SUM[20]) );
  AOI21X1 U647 ( .A0(n162), .A1(n158), .B0(n159), .Y(n157) );
  XOR2X1 U648 ( .A(n144), .B(n18), .Y(SUM[22]) );
  XNOR2X1 U649 ( .A(n130), .B(n16), .Y(SUM[24]) );
  NAND2X1 U650 ( .A(n277), .B(n129), .Y(n16) );
  OAI21XL U651 ( .A0(n144), .A1(n131), .B0(n132), .Y(n130) );
  NAND2X1 U652 ( .A(n428), .B(n151), .Y(n19) );
endmodule


module CONV ( clk, reset, busy, ready, iaddr, idata, cwr, caddr_wr, cdata_wr, 
        crd, caddr_rd, cdata_rd, csel );
  output [11:0] iaddr;
  input [19:0] idata;
  output [11:0] caddr_wr;
  output [19:0] cdata_wr;
  output [11:0] caddr_rd;
  input [19:0] cdata_rd;
  output [2:0] csel;
  input clk, reset, ready;
  output busy, cwr, crd;
  wire   n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N157, N158, N159, N160, N161, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N365, N366, N367, N368, N369, N370, N371, N372, N373,
         N374, N375, N424, N425, N426, N427, N428, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N609, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N681,
         N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692,
         N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704,
         N705, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744,
         N745, N937, N938, N939, N940, n51, n52, n55, n68, n69, n70, n71, n72,
         n76, n77, n78, n79, n80, n81, n82, n104, n106, n107, n108, n109, n110,
         n111, n112, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, \mul[9] , \mul[8] , \mul[7] , \mul[6] ,
         \mul[5] , \mul[4] , \mul[3] , \mul[39] , \mul[38] , \mul[37] ,
         \mul[36] , \mul[35] , \mul[34] , \mul[33] , \mul[32] , \mul[31] ,
         \mul[30] , \mul[2] , \mul[29] , \mul[28] , \mul[27] , \mul[26] ,
         \mul[25] , \mul[24] , \mul[23] , \mul[22] , \mul[21] , \mul[20] ,
         \mul[1] , \mul[19] , \mul[18] , \mul[17] , \mul[16] , \mul[15] ,
         \mul[14] , \mul[13] , \mul[12] , \mul[11] , \mul[10] , \mul[0] ,
         \sub_172/carry[7] , \sub_172/carry[8] , \sub_172/carry[9] ,
         \sub_172/carry[10] , \sub_172/carry[11] , \add_153/carry[2] ,
         \add_153/carry[3] , \add_153/carry[4] , \add_153/carry[5] ,
         \add_153/carry[6] , \add_103/carry[7] , \add_90/carry[2] ,
         \add_90/carry[3] , \add_90/carry[4] , \add_90/carry[5] ,
         \add_90/carry[6] , \sub_62/carry[7] , \sub_62/carry[8] ,
         \sub_62/carry[9] , \sub_62/carry[10] , \sub_62/carry[11] ,
         \sub_57/carry[11] , \sub_57/carry[10] , \sub_57/carry[9] ,
         \sub_57/carry[8] , \sub_54/carry[2] , \sub_54/carry[3] ,
         \sub_54/carry[4] , \sub_54/carry[5] , \sub_54/carry[6] ,
         \sub_54/carry[8] , \sub_54/carry[9] , \sub_54/carry[10] ,
         \sub_54/carry[11] , \r406/carry[4] , \r406/carry[3] , \r406/carry[2] ,
         n538, n539, n540, n541, n561, n563, n571, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n671, n673, n675, n677, n679, n681,
         n683, n685, n687, n689, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104;
  wire   [19:0] data;
  wire   [19:0] kernel;
  wire   [4:0] state;
  wire   [39:0] sum;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign csel[2] = 1'b0;

  CONV_DW01_dec_0 sub_69 ( .A({n692, n671, n673, n675, n677, n679, n681, n683, 
        n685, n687, n689, caddr_wr[0]}), .SUM({N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219, N218, N217}) );
  CONV_DW_cmp_4 r400 ( .A(cdata_rd), .B({n1126, n1127, n1128, n1129, n1130, 
        n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
        n1141, n1142, n1143, n1144, n1145}), .TC(1'b0), .GE_LT(1'b0), 
        .GE_GT_EQ(1'b1), .GE_LT_GT_LE(N705) );
  CONV_DW01_inc_1 r398 ( .A({n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
        n1154, n1155, n1156, n1157, n1158}), .SUM({N692, N691, N690, N689, 
        N688, N687, N686, N685, N684, N683, N682, N681}) );
  CONV_DW01_inc_2 r392 ( .A({n692, n671, n673, n675, n677, n679, n681, n683, 
        n685, n687, n689, caddr_wr[0]}), .SUM({N323, N322, N321, N320, N319, 
        N318, N317, N316, N315, N314, N313, SYNOPSYS_UNCONNECTED__0}) );
  CONV_DW_mult_tc_2 mult_27 ( .a(data), .b(kernel), .product({\mul[39] , 
        \mul[38] , \mul[37] , \mul[36] , \mul[35] , \mul[34] , \mul[33] , 
        \mul[32] , \mul[31] , \mul[30] , \mul[29] , \mul[28] , \mul[27] , 
        \mul[26] , \mul[25] , \mul[24] , \mul[23] , \mul[22] , \mul[21] , 
        \mul[20] , \mul[19] , \mul[18] , \mul[17] , \mul[16] , \mul[15] , 
        \mul[14] , \mul[13] , \mul[12] , \mul[11] , \mul[10] , \mul[9] , 
        \mul[8] , \mul[7] , \mul[6] , \mul[5] , \mul[4] , \mul[3] , \mul[2] , 
        \mul[1] , \mul[0] }) );
  CONV_DW01_add_8 r390 ( .A({sum[39:20], N631, N630, N629, N628, sum[15:0]}), 
        .B({\mul[39] , \mul[38] , \mul[37] , \mul[36] , \mul[35] , \mul[34] , 
        \mul[33] , \mul[32] , \mul[31] , \mul[30] , \mul[29] , \mul[28] , 
        \mul[27] , \mul[26] , \mul[25] , \mul[24] , \mul[23] , \mul[22] , 
        \mul[21] , \mul[20] , \mul[19] , \mul[18] , \mul[17] , \mul[16] , 
        \mul[15] , \mul[14] , \mul[13] , \mul[12] , \mul[11] , \mul[10] , 
        \mul[9] , \mul[8] , \mul[7] , \mul[6] , \mul[5] , \mul[4] , \mul[3] , 
        \mul[2] , \mul[1] , \mul[0] }), .CI(1'b0), .SUM({N215, N214, N213, 
        N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, 
        N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, 
        N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, 
        N176}) );
  DFFRX1 \sum_reg[39]  ( .D(n467), .CK(clk), .RN(n705), .Q(sum[39]), .QN(n1096) );
  DFFRX1 \sum_reg[38]  ( .D(n466), .CK(clk), .RN(n705), .Q(sum[38]), .QN(n1095) );
  DFFRX2 \sum_reg[27]  ( .D(n455), .CK(clk), .RN(n714), .Q(sum[27]), .QN(n1084) );
  DFFRX2 \sum_reg[31]  ( .D(n459), .CK(clk), .RN(n714), .Q(sum[31]), .QN(n1088) );
  DFFRX2 \sum_reg[29]  ( .D(n457), .CK(clk), .RN(n714), .Q(sum[29]), .QN(n1086) );
  DFFRX1 \sum_reg[14]  ( .D(n422), .CK(clk), .RN(n713), .Q(sum[14]), .QN(n1053) );
  DFFRX1 \sum_reg[13]  ( .D(n421), .CK(clk), .RN(n713), .Q(sum[13]), .QN(n1052) );
  DFFRX1 \sum_reg[12]  ( .D(n420), .CK(clk), .RN(n713), .Q(sum[12]), .QN(n1051) );
  DFFRX1 \sum_reg[11]  ( .D(n419), .CK(clk), .RN(n713), .Q(sum[11]), .QN(n1050) );
  DFFRX1 \sum_reg[10]  ( .D(n418), .CK(clk), .RN(n713), .Q(sum[10]), .QN(n1049) );
  DFFRX1 \sum_reg[9]  ( .D(n417), .CK(clk), .RN(n712), .Q(sum[9]), .QN(n1048)
         );
  DFFRX1 \sum_reg[7]  ( .D(n415), .CK(clk), .RN(n712), .Q(sum[7]), .QN(n1046)
         );
  DFFRX2 \sum_reg[23]  ( .D(n451), .CK(clk), .RN(n714), .Q(sum[23]), .QN(n1080) );
  DFFRX1 \caddr_wr_reg[6]  ( .D(n504), .CK(clk), .RN(n703), .Q(n1125), .QN(n72) );
  DFFRX1 \caddr_wr_reg[8]  ( .D(n502), .CK(clk), .RN(n703), .Q(n1123), .QN(n70) );
  DFFRX1 \caddr_wr_reg[7]  ( .D(n503), .CK(clk), .RN(n703), .Q(n1124), .QN(n71) );
  DFFRX1 \caddr_wr_reg[9]  ( .D(n501), .CK(clk), .RN(n703), .Q(n1122), .QN(n69) );
  DFFRX1 \sum_reg[8]  ( .D(n416), .CK(clk), .RN(n712), .Q(sum[8]), .QN(n1047)
         );
  DFFRX1 \sum_reg[6]  ( .D(n414), .CK(clk), .RN(n712), .Q(sum[6]), .QN(n1045)
         );
  DFFRX1 \sum_reg[5]  ( .D(n413), .CK(clk), .RN(n712), .Q(sum[5]), .QN(n1044)
         );
  DFFRX1 \sum_reg[4]  ( .D(n412), .CK(clk), .RN(n712), .Q(sum[4]), .QN(n1043)
         );
  DFFRX1 \sum_reg[3]  ( .D(n411), .CK(clk), .RN(n712), .Q(sum[3]), .QN(n1042)
         );
  DFFRX1 \sum_reg[2]  ( .D(n410), .CK(clk), .RN(n712), .Q(sum[2]), .QN(n1041)
         );
  DFFRX1 \sum_reg[1]  ( .D(n409), .CK(clk), .RN(n712), .Q(sum[1]), .QN(n1040)
         );
  DFFRX1 \caddr_wr_reg[11]  ( .D(n511), .CK(clk), .RN(n703), .Q(n1120), .QN(
        n55) );
  DFFRX1 \caddr_wr_reg[10]  ( .D(n500), .CK(clk), .RN(n704), .Q(n1121), .QN(
        n68) );
  DFFRX2 \sum_reg[21]  ( .D(n449), .CK(clk), .RN(n713), .Q(sum[21]), .QN(n1078) );
  DFFRX1 \caddr_wr_reg[4]  ( .D(n506), .CK(clk), .RN(n703), .Q(N154), .QN(n77)
         );
  DFFRX1 \caddr_wr_reg[5]  ( .D(n505), .CK(clk), .RN(n703), .Q(N155), .QN(n76)
         );
  DFFRX1 \sum_reg[0]  ( .D(n408), .CK(clk), .RN(n712), .Q(sum[0]), .QN(n1039)
         );
  DFFRX1 \caddr_wr_reg[2]  ( .D(n508), .CK(clk), .RN(n703), .Q(N152), .QN(n79)
         );
  DFFRX1 \caddr_wr_reg[3]  ( .D(n507), .CK(clk), .RN(n703), .Q(N153), .QN(n78)
         );
  DFFRX1 \kernel_reg[19]  ( .D(n512), .CK(clk), .RN(n710), .Q(kernel[19]), 
        .QN(n1019) );
  DFFRX1 \kernel_reg[18]  ( .D(n513), .CK(clk), .RN(n710), .Q(kernel[18]), 
        .QN(n1020) );
  DFFRX1 \caddr_wr_reg[0]  ( .D(n510), .CK(clk), .RN(n703), .Q(N150), .QN(n81)
         );
  DFFRX1 \caddr_wr_reg[1]  ( .D(n509), .CK(clk), .RN(n703), .Q(N151), .QN(n80)
         );
  ADDHXL \r406/U1_1_3  ( .A(state[3]), .B(\r406/carry[3] ), .CO(
        \r406/carry[4] ), .S(N939) );
  ADDHXL \r406/U1_1_2  ( .A(state[2]), .B(\r406/carry[2] ), .CO(
        \r406/carry[3] ), .S(N938) );
  ADDHXL \r406/U1_1_1  ( .A(state[1]), .B(state[0]), .CO(\r406/carry[2] ), .S(
        N937) );
  DFFRX1 \sum_reg[32]  ( .D(n460), .CK(clk), .RN(n714), .Q(sum[32]), .QN(n1089) );
  DFFRX1 \sum_reg[30]  ( .D(n458), .CK(clk), .RN(n714), .Q(sum[30]), .QN(n1087) );
  DFFRX1 \sum_reg[22]  ( .D(n450), .CK(clk), .RN(n714), .Q(sum[22]), .QN(n1079) );
  DFFRX1 \sum_reg[25]  ( .D(n453), .CK(clk), .RN(n714), .Q(sum[25]), .QN(n1082) );
  DFFRX1 \sum_reg[19]  ( .D(n447), .CK(clk), .RN(n713), .Q(N631), .QN(n1076)
         );
  DFFRX1 \sum_reg[17]  ( .D(n445), .CK(clk), .RN(n713), .Q(N629), .QN(n1074)
         );
  DFFRX2 \kernel_reg[16]  ( .D(n515), .CK(clk), .RN(n710), .Q(kernel[16]), 
        .QN(n1022) );
  DFFRX2 \kernel_reg[14]  ( .D(n517), .CK(clk), .RN(n710), .Q(kernel[14]), 
        .QN(n1023) );
  DFFRX2 \kernel_reg[12]  ( .D(n519), .CK(clk), .RN(n709), .Q(kernel[12]), 
        .QN(n1024) );
  DFFRX2 \kernel_reg[8]  ( .D(n523), .CK(clk), .RN(n709), .Q(kernel[8]), .QN(
        n1026) );
  DFFRX2 \kernel_reg[6]  ( .D(n525), .CK(clk), .RN(n709), .Q(kernel[6]), .QN(
        n52) );
  DFFRX2 \kernel_reg[7]  ( .D(n524), .CK(clk), .RN(n709), .Q(kernel[7]), .QN(
        n1027) );
  DFFRX2 \kernel_reg[3]  ( .D(n528), .CK(clk), .RN(n709), .Q(kernel[3]), .QN(
        n1030) );
  DFFRX4 \data_reg[19]  ( .D(n487), .CK(clk), .RN(n712), .Q(data[19]) );
  DFFRX4 \data_reg[15]  ( .D(n483), .CK(clk), .RN(n711), .Q(data[15]) );
  DFFRX4 \data_reg[10]  ( .D(n478), .CK(clk), .RN(n711), .Q(data[10]) );
  DFFRX4 \data_reg[6]  ( .D(n474), .CK(clk), .RN(n711), .Q(data[6]) );
  DFFRX4 \data_reg[9]  ( .D(n477), .CK(clk), .RN(n711), .Q(data[9]) );
  DFFRX4 \data_reg[7]  ( .D(n475), .CK(clk), .RN(n711), .Q(data[7]) );
  DFFRX4 \data_reg[5]  ( .D(n473), .CK(clk), .RN(n710), .Q(data[5]) );
  DFFRX1 \sum_reg[36]  ( .D(n464), .CK(clk), .RN(n705), .Q(sum[36]), .QN(n1093) );
  DFFRX1 \sum_reg[28]  ( .D(n456), .CK(clk), .RN(n714), .Q(sum[28]), .QN(n1085) );
  DFFRX1 \sum_reg[26]  ( .D(n454), .CK(clk), .RN(n714), .Q(sum[26]), .QN(n1083) );
  DFFRX1 \sum_reg[33]  ( .D(n461), .CK(clk), .RN(n714), .Q(sum[33]), .QN(n1090) );
  DFFRX1 \sum_reg[18]  ( .D(n446), .CK(clk), .RN(n713), .Q(N630), .QN(n1075)
         );
  DFFRX1 \sum_reg[37]  ( .D(n465), .CK(clk), .RN(n705), .Q(sum[37]), .QN(n1094) );
  DFFRX1 \sum_reg[35]  ( .D(n463), .CK(clk), .RN(n708), .Q(sum[35]), .QN(n1092) );
  DFFRX1 \sum_reg[24]  ( .D(n452), .CK(clk), .RN(n714), .Q(sum[24]), .QN(n1081) );
  DFFRX1 \caddr_rd_reg[10]  ( .D(n397), .CK(clk), .RN(n707), .Q(n1148), .QN(
        n1035) );
  DFFRX1 \caddr_rd_reg[2]  ( .D(n405), .CK(clk), .RN(n707), .Q(n1156), .QN(
        n110) );
  DFFRX1 \caddr_rd_reg[3]  ( .D(n404), .CK(clk), .RN(n707), .Q(n1155), .QN(
        n109) );
  DFFRX1 \caddr_rd_reg[4]  ( .D(n403), .CK(clk), .RN(n707), .Q(n1154), .QN(
        n108) );
  DFFRX1 \caddr_rd_reg[5]  ( .D(n402), .CK(clk), .RN(n708), .Q(n1153), .QN(
        n107) );
  DFFRX1 \caddr_rd_reg[6]  ( .D(n401), .CK(clk), .RN(n708), .Q(n1152), .QN(
        n106) );
  DFFRX1 \caddr_rd_reg[9]  ( .D(n398), .CK(clk), .RN(n708), .Q(n1149), .QN(
        n1036) );
  DFFRX1 \caddr_rd_reg[7]  ( .D(n400), .CK(clk), .RN(n708), .Q(n1151), .QN(
        n1038) );
  DFFRX1 \caddr_rd_reg[8]  ( .D(n399), .CK(clk), .RN(n708), .Q(n1150), .QN(
        n1037) );
  DFFRX2 \cdata_wr_reg[12]  ( .D(n429), .CK(clk), .RN(n706), .Q(n1133), .QN(
        n1060) );
  DFFRX2 \cdata_wr_reg[19]  ( .D(n442), .CK(clk), .RN(n705), .Q(n1126), .QN(
        n104) );
  DFFRX2 \cdata_wr_reg[17]  ( .D(n424), .CK(clk), .RN(n705), .Q(n1128), .QN(
        n1055) );
  DFFRX2 \cdata_wr_reg[14]  ( .D(n427), .CK(clk), .RN(n706), .Q(n1131), .QN(
        n1058) );
  DFFRX2 \cdata_wr_reg[8]  ( .D(n433), .CK(clk), .RN(n706), .Q(n1137), .QN(
        n1064) );
  DFFRX2 \cdata_wr_reg[5]  ( .D(n436), .CK(clk), .RN(n706), .Q(n1140), .QN(
        n1067) );
  DFFRX2 \cdata_wr_reg[3]  ( .D(n438), .CK(clk), .RN(n707), .Q(n1142), .QN(
        n1069) );
  DFFRX1 \caddr_rd_reg[11]  ( .D(n396), .CK(clk), .RN(n707), .Q(n1147), .QN(
        n1034) );
  DFFRX2 \cdata_wr_reg[18]  ( .D(n423), .CK(clk), .RN(n705), .Q(n1127), .QN(
        n1054) );
  DFFRX2 \cdata_wr_reg[0]  ( .D(n441), .CK(clk), .RN(n707), .Q(n1145), .QN(
        n1072) );
  DFFRX2 \cdata_wr_reg[13]  ( .D(n428), .CK(clk), .RN(n706), .Q(n1132), .QN(
        n1059) );
  DFFRX1 \iaddr_reg[0]  ( .D(n499), .CK(clk), .RN(n704), .Q(n1118), .QN(n571)
         );
  DFFRX2 \cdata_wr_reg[11]  ( .D(n430), .CK(clk), .RN(n706), .Q(n1134), .QN(
        n1061) );
  DFFRX2 \cdata_wr_reg[15]  ( .D(n426), .CK(clk), .RN(n706), .Q(n1130), .QN(
        n1057) );
  DFFRX2 \cdata_wr_reg[9]  ( .D(n432), .CK(clk), .RN(n706), .Q(n1136), .QN(
        n1063) );
  DFFRX2 \cdata_wr_reg[1]  ( .D(n440), .CK(clk), .RN(n707), .Q(n1144), .QN(
        n1071) );
  DFFRX2 \cdata_wr_reg[6]  ( .D(n435), .CK(clk), .RN(n706), .Q(n1139), .QN(
        n1066) );
  DFFRX1 cwr_reg ( .D(n392), .CK(clk), .RN(n708), .Q(n1119), .QN(n563) );
  DFFRX1 \csel_reg[0]  ( .D(n394), .CK(clk), .RN(n708), .Q(n1160), .QN(n561)
         );
  DFFRX1 \csel_reg[1]  ( .D(n395), .CK(clk), .RN(n708), .Q(n1159), .QN(n1033)
         );
  DFFRX1 \iaddr_reg[8]  ( .D(n491), .CK(clk), .RN(n705), .Q(n1110), .QN(n1100)
         );
  DFFRX1 \iaddr_reg[9]  ( .D(n490), .CK(clk), .RN(n704), .Q(n1109), .QN(n1099)
         );
  DFFRX1 \iaddr_reg[10]  ( .D(n489), .CK(clk), .RN(n704), .Q(n1108), .QN(n1098) );
  DFFRX1 \iaddr_reg[11]  ( .D(n488), .CK(clk), .RN(n704), .Q(n1107), .QN(n1097) );
  DFFRX1 \iaddr_reg[4]  ( .D(n495), .CK(clk), .RN(n705), .Q(n1114), .QN(n1104)
         );
  DFFRX1 \iaddr_reg[5]  ( .D(n494), .CK(clk), .RN(n705), .Q(n1113), .QN(n1103)
         );
  DFFRX1 \iaddr_reg[6]  ( .D(n493), .CK(clk), .RN(n705), .Q(n1112), .QN(n1102)
         );
  DFFRX1 \iaddr_reg[7]  ( .D(n492), .CK(clk), .RN(n705), .Q(n1111), .QN(n1101)
         );
  DFFRX1 \iaddr_reg[1]  ( .D(n498), .CK(clk), .RN(n704), .Q(n1117), .QN(n1018)
         );
  DFFRX1 \iaddr_reg[2]  ( .D(n497), .CK(clk), .RN(n704), .Q(n1116), .QN(n1017)
         );
  DFFRX1 \iaddr_reg[3]  ( .D(n496), .CK(clk), .RN(n704), .Q(n1115), .QN(n1016)
         );
  DFFRX1 crd_reg ( .D(n393), .CK(clk), .RN(n708), .Q(n1146), .QN(n1032) );
  DFFRX1 \caddr_rd_reg[1]  ( .D(n406), .CK(clk), .RN(n707), .Q(n1157), .QN(
        n111) );
  DFFRX2 \cdata_wr_reg[10]  ( .D(n431), .CK(clk), .RN(n706), .Q(n1135), .QN(
        n1062) );
  DFFRX2 \cdata_wr_reg[16]  ( .D(n425), .CK(clk), .RN(n706), .Q(n1129), .QN(
        n1056) );
  DFFRX1 \state_reg[0]  ( .D(n537), .CK(clk), .RN(n777), .Q(state[0]), .QN(
        n783) );
  DFFRX1 \state_reg[4]  ( .D(n536), .CK(clk), .RN(n777), .Q(state[4]), .QN(
        n788) );
  DFFRX1 \state_reg[1]  ( .D(n534), .CK(clk), .RN(n777), .Q(state[1]), .QN(
        n1015) );
  DFFRX1 \state_reg[2]  ( .D(n533), .CK(clk), .RN(n777), .Q(state[2]), .QN(
        n797) );
  DFFRX1 \data_reg[0]  ( .D(n468), .CK(clk), .RN(n777), .Q(data[0]) );
  DFFRX1 \sum_reg[15]  ( .D(n443), .CK(clk), .RN(n777), .Q(sum[15]), .QN(n746)
         );
  DFFSRX1 \state_reg[3]  ( .D(n532), .CK(clk), .SN(1'b1), .RN(n777), .Q(
        state[3]), .QN(n799) );
  DFFRX2 busy_reg ( .D(n535), .CK(clk), .RN(n777), .Q(n1106), .QN(n82) );
  DFFRX1 \sum_reg[16]  ( .D(n444), .CK(clk), .RN(n713), .Q(N628), .QN(n1073)
         );
  DFFRX1 \kernel_reg[13]  ( .D(n518), .CK(clk), .RN(n709), .Q(kernel[13]), 
        .QN(n541) );
  DFFRX1 \kernel_reg[1]  ( .D(n530), .CK(clk), .RN(n708), .Q(kernel[1]), .QN(
        n540) );
  DFFRX1 \kernel_reg[9]  ( .D(n522), .CK(clk), .RN(n709), .Q(kernel[9]), .QN(
        n539) );
  DFFRX1 \caddr_rd_reg[0]  ( .D(n407), .CK(clk), .RN(n707), .Q(n1158), .QN(
        n112) );
  DFFRX1 \sum_reg[20]  ( .D(n448), .CK(clk), .RN(n713), .Q(sum[20]), .QN(n1077) );
  DFFRX2 \data_reg[1]  ( .D(n469), .CK(clk), .RN(n710), .Q(data[1]) );
  DFFRX2 \cdata_wr_reg[7]  ( .D(n434), .CK(clk), .RN(n706), .Q(n1138), .QN(
        n1065) );
  DFFRX1 \kernel_reg[15]  ( .D(n516), .CK(clk), .RN(n710), .Q(kernel[15]), 
        .QN(n51) );
  DFFRX1 \kernel_reg[10]  ( .D(n521), .CK(clk), .RN(n709), .Q(kernel[10]), 
        .QN(n1025) );
  DFFRX2 \data_reg[14]  ( .D(n482), .CK(clk), .RN(n711), .Q(data[14]) );
  DFFRX2 \data_reg[18]  ( .D(n486), .CK(clk), .RN(n712), .Q(data[18]) );
  DFFRX2 \data_reg[16]  ( .D(n484), .CK(clk), .RN(n711), .Q(data[16]) );
  DFFRX2 \data_reg[17]  ( .D(n485), .CK(clk), .RN(n711), .Q(data[17]) );
  DFFRX2 \kernel_reg[5]  ( .D(n526), .CK(clk), .RN(n709), .Q(kernel[5]), .QN(
        n1028) );
  DFFRX1 \kernel_reg[0]  ( .D(n531), .CK(clk), .RN(n708), .Q(kernel[0]), .QN(
        n1031) );
  DFFRX2 \kernel_reg[2]  ( .D(n529), .CK(clk), .RN(n709), .Q(kernel[2]) );
  DFFRX2 \kernel_reg[11]  ( .D(n520), .CK(clk), .RN(n709), .Q(kernel[11]) );
  DFFRX2 \data_reg[12]  ( .D(n480), .CK(clk), .RN(n711), .Q(data[12]) );
  DFFRX2 \data_reg[8]  ( .D(n476), .CK(clk), .RN(n711), .Q(data[8]) );
  DFFRX2 \data_reg[2]  ( .D(n470), .CK(clk), .RN(n710), .Q(data[2]) );
  DFFRX2 \data_reg[4]  ( .D(n472), .CK(clk), .RN(n710), .Q(data[4]) );
  DFFRX2 \data_reg[13]  ( .D(n481), .CK(clk), .RN(n711), .Q(data[13]) );
  DFFRX2 \data_reg[11]  ( .D(n479), .CK(clk), .RN(n711), .Q(data[11]) );
  DFFRX2 \data_reg[3]  ( .D(n471), .CK(clk), .RN(n710), .Q(data[3]) );
  DFFRX2 \kernel_reg[17]  ( .D(n514), .CK(clk), .RN(n710), .Q(kernel[17]), 
        .QN(n1021) );
  DFFRX2 \kernel_reg[4]  ( .D(n527), .CK(clk), .RN(n709), .Q(kernel[4]), .QN(
        n1029) );
  DFFRX1 \sum_reg[34]  ( .D(n462), .CK(clk), .RN(n702), .Q(sum[34]), .QN(n1091) );
  DFFRX1 \cdata_wr_reg[4]  ( .D(n437), .CK(clk), .RN(n707), .Q(n1141), .QN(
        n1068) );
  DFFRX1 \cdata_wr_reg[2]  ( .D(n439), .CK(clk), .RN(n707), .Q(n1143), .QN(
        n1070) );
  OAI2BB2X1 U482 ( .B0(n1094), .B1(n774), .A0N(N213), .A1N(n773), .Y(n465) );
  OAI31XL U483 ( .A0(n720), .A1(n719), .A2(n718), .B0(n1106), .Y(n723) );
  BUFX12 U484 ( .A(n776), .Y(n653) );
  BUFX4 U485 ( .A(n907), .Y(n666) );
  OAI2BB2XL U486 ( .B0(n1091), .B1(n699), .A0N(N210), .A1N(n697), .Y(n462) );
  OAI2BB2XL U487 ( .B0(n1090), .B1(n699), .A0N(N209), .A1N(n696), .Y(n461) );
  AOI2BB1X1 U488 ( .A0N(n1031), .A1N(n695), .B0(n597), .Y(n741) );
  OAI2BB2XL U489 ( .B0(n1089), .B1(n699), .A0N(N208), .A1N(n697), .Y(n460) );
  OAI2BB2XL U490 ( .B0(n1088), .B1(n698), .A0N(N207), .A1N(n697), .Y(n459) );
  AND2X2 U491 ( .A(n962), .B(state[3]), .Y(n538) );
  INVX3 U492 ( .A(reset), .Y(n777) );
  NAND2XL U494 ( .A(cdata_rd[2]), .B(n666), .Y(n912) );
  INVX12 U495 ( .A(n1065), .Y(cdata_wr[7]) );
  INVX12 U496 ( .A(n1056), .Y(cdata_wr[16]) );
  INVX12 U497 ( .A(n1070), .Y(cdata_wr[2]) );
  INVX12 U498 ( .A(n1062), .Y(cdata_wr[10]) );
  BUFX12 U499 ( .A(n1157), .Y(caddr_rd[1]) );
  BUFX12 U500 ( .A(n1146), .Y(crd) );
  BUFX12 U501 ( .A(n1115), .Y(iaddr[3]) );
  BUFX12 U502 ( .A(n1116), .Y(iaddr[2]) );
  BUFX12 U503 ( .A(n1117), .Y(iaddr[1]) );
  BUFX12 U504 ( .A(n1111), .Y(iaddr[7]) );
  BUFX12 U505 ( .A(n1112), .Y(iaddr[6]) );
  BUFX12 U506 ( .A(n1113), .Y(iaddr[5]) );
  BUFX12 U507 ( .A(n1114), .Y(iaddr[4]) );
  BUFX12 U508 ( .A(n1107), .Y(iaddr[11]) );
  BUFX12 U509 ( .A(n1108), .Y(iaddr[10]) );
  BUFX12 U510 ( .A(n1109), .Y(iaddr[9]) );
  BUFX12 U511 ( .A(n1110), .Y(iaddr[8]) );
  BUFX12 U512 ( .A(n1159), .Y(csel[1]) );
  NOR2X2 U513 ( .A(state[0]), .B(state[1]), .Y(n808) );
  INVX12 U514 ( .A(n561), .Y(csel[0]) );
  INVX12 U515 ( .A(n563), .Y(cwr) );
  INVX12 U516 ( .A(n1066), .Y(cdata_wr[6]) );
  INVX12 U517 ( .A(n1071), .Y(cdata_wr[1]) );
  INVX12 U518 ( .A(n1068), .Y(cdata_wr[4]) );
  INVX12 U519 ( .A(n1063), .Y(cdata_wr[9]) );
  INVX12 U520 ( .A(n1057), .Y(cdata_wr[15]) );
  INVX12 U521 ( .A(n1061), .Y(cdata_wr[11]) );
  INVX12 U522 ( .A(n571), .Y(iaddr[0]) );
  INVX12 U523 ( .A(n1059), .Y(cdata_wr[13]) );
  INVX12 U524 ( .A(n1072), .Y(cdata_wr[0]) );
  INVX12 U525 ( .A(n1054), .Y(cdata_wr[18]) );
  BUFX12 U526 ( .A(n1147), .Y(caddr_rd[11]) );
  INVX12 U527 ( .A(n1069), .Y(cdata_wr[3]) );
  INVX12 U528 ( .A(n1067), .Y(cdata_wr[5]) );
  INVX12 U529 ( .A(n1064), .Y(cdata_wr[8]) );
  INVX12 U530 ( .A(n1058), .Y(cdata_wr[14]) );
  INVX12 U531 ( .A(n1055), .Y(cdata_wr[17]) );
  INVX12 U532 ( .A(n104), .Y(cdata_wr[19]) );
  INVX12 U533 ( .A(n1060), .Y(cdata_wr[12]) );
  BUFX12 U534 ( .A(n1150), .Y(caddr_rd[8]) );
  BUFX12 U535 ( .A(n1151), .Y(caddr_rd[7]) );
  BUFX12 U536 ( .A(n1149), .Y(caddr_rd[9]) );
  BUFX12 U537 ( .A(n1152), .Y(caddr_rd[6]) );
  BUFX12 U538 ( .A(n1153), .Y(caddr_rd[5]) );
  BUFX12 U539 ( .A(n1154), .Y(caddr_rd[4]) );
  BUFX12 U540 ( .A(n1155), .Y(caddr_rd[3]) );
  BUFX12 U541 ( .A(n1156), .Y(caddr_rd[2]) );
  BUFX12 U542 ( .A(n1148), .Y(caddr_rd[10]) );
  INVX12 U543 ( .A(n112), .Y(caddr_rd[0]) );
  NAND2XL U544 ( .A(n538), .B(n806), .Y(n946) );
  NAND2XL U545 ( .A(n902), .B(n806), .Y(n897) );
  NAND2XL U546 ( .A(n956), .B(n806), .Y(n895) );
  NAND2XL U547 ( .A(n1003), .B(n806), .Y(n953) );
  NAND2XL U548 ( .A(n902), .B(n808), .Y(n894) );
  OAI2BB2XL U549 ( .B0(n1092), .B1(n774), .A0N(N211), .A1N(n696), .Y(n463) );
  OAI2BB2XL U550 ( .B0(n1085), .B1(n698), .A0N(N204), .A1N(n697), .Y(n456) );
  AOI211XL U551 ( .A0(n665), .A1(n1118), .B0(n838), .C0(n839), .Y(n836) );
  NAND2XL U552 ( .A(n1148), .B(n630), .Y(n649) );
  NAND2BXL U553 ( .AN(n1158), .B(n973), .Y(n969) );
  OR2XL U554 ( .A(n1153), .B(\add_153/carry[5] ), .Y(\add_153/carry[6] ) );
  OR2XL U555 ( .A(n1157), .B(n1158), .Y(\add_153/carry[2] ) );
  OR2XL U556 ( .A(n1156), .B(\add_153/carry[2] ), .Y(\add_153/carry[3] ) );
  OR2XL U557 ( .A(n1155), .B(\add_153/carry[3] ), .Y(\add_153/carry[4] ) );
  OR2XL U558 ( .A(n1154), .B(\add_153/carry[4] ), .Y(\add_153/carry[5] ) );
  OR2XL U559 ( .A(n1150), .B(\sub_172/carry[8] ), .Y(\sub_172/carry[9] ) );
  OR2XL U560 ( .A(n1151), .B(\sub_172/carry[7] ), .Y(\sub_172/carry[8] ) );
  OR2XL U561 ( .A(n1152), .B(n625), .Y(\sub_172/carry[7] ) );
  OR2XL U562 ( .A(n1149), .B(\sub_172/carry[9] ), .Y(\sub_172/carry[10] ) );
  OR2XL U563 ( .A(n1148), .B(\sub_172/carry[10] ), .Y(\sub_172/carry[11] ) );
  AND2XL U564 ( .A(n1157), .B(n1158), .Y(n634) );
  AND2XL U565 ( .A(n1149), .B(n629), .Y(n630) );
  AND2XL U566 ( .A(n1152), .B(\add_153/carry[6] ), .Y(n627) );
  AND2XL U567 ( .A(n1151), .B(n627), .Y(n628) );
  AND2XL U568 ( .A(n1150), .B(n628), .Y(n629) );
  AND2XL U569 ( .A(n1154), .B(n632), .Y(n631) );
  AND2XL U570 ( .A(n1155), .B(n633), .Y(n632) );
  AND2XL U571 ( .A(n1156), .B(n634), .Y(n633) );
  AND2XL U572 ( .A(n1153), .B(n631), .Y(n625) );
  MXI2XL U573 ( .A(n1119), .B(n833), .S0(n1006), .Y(n1013) );
  MXI2XL U574 ( .A(n1160), .B(n952), .S0(n1006), .Y(n1008) );
  NOR2XL U575 ( .A(n785), .B(n787), .Y(n791) );
  MXI2XL U576 ( .A(n806), .B(n807), .S0(state[2]), .Y(n805) );
  MXI2XL U577 ( .A(n1010), .B(n1032), .S0(n1011), .Y(n393) );
  NAND2XL U578 ( .A(n785), .B(n794), .Y(n793) );
  CLKBUFX3 U579 ( .A(n740), .Y(n694) );
  BUFX20 U580 ( .A(n775), .Y(n654) );
  CLKINVX4 U581 ( .A(n753), .Y(n775) );
  CLKINVX4 U582 ( .A(n754), .Y(n776) );
  CLKINVX1 U583 ( .A(n731), .Y(n740) );
  CLKINVX1 U584 ( .A(n723), .Y(n774) );
  CLKBUFX3 U585 ( .A(n837), .Y(n665) );
  CLKINVX1 U586 ( .A(n722), .Y(n773) );
  OAI2BB2X1 U587 ( .B0(n1096), .B1(n699), .A0N(N215), .A1N(n696), .Y(n467) );
  AOI221X2 U588 ( .A0(n949), .A1(n950), .B0(n833), .B1(n104), .C0(n82), .Y(
        n904) );
  BUFX20 U589 ( .A(n904), .Y(n667) );
  NAND2XL U590 ( .A(n731), .B(kernel[11]), .Y(n728) );
  MXI2XL U591 ( .A(kernel[2]), .B(n809), .S0(n693), .Y(n626) );
  MX2XL U592 ( .A(data[0]), .B(idata[0]), .S0(n693), .Y(n468) );
  MX2XL U593 ( .A(data[1]), .B(idata[1]), .S0(n693), .Y(n469) );
  MX2XL U594 ( .A(data[2]), .B(idata[2]), .S0(n693), .Y(n470) );
  MX2XL U595 ( .A(data[3]), .B(idata[3]), .S0(n693), .Y(n471) );
  MX2XL U596 ( .A(data[19]), .B(idata[19]), .S0(n693), .Y(n487) );
  MX2XL U597 ( .A(data[4]), .B(idata[4]), .S0(n694), .Y(n472) );
  MX2XL U598 ( .A(data[5]), .B(idata[5]), .S0(n694), .Y(n473) );
  MX2XL U599 ( .A(data[6]), .B(idata[6]), .S0(n694), .Y(n474) );
  MX2XL U600 ( .A(data[7]), .B(idata[7]), .S0(n694), .Y(n475) );
  MX2XL U601 ( .A(data[8]), .B(idata[8]), .S0(n694), .Y(n476) );
  MX2XL U602 ( .A(data[9]), .B(idata[9]), .S0(n694), .Y(n477) );
  MX2XL U603 ( .A(data[10]), .B(idata[10]), .S0(n694), .Y(n478) );
  MX2XL U604 ( .A(data[11]), .B(idata[11]), .S0(n694), .Y(n479) );
  MX2XL U605 ( .A(data[12]), .B(idata[12]), .S0(n694), .Y(n480) );
  MX2XL U606 ( .A(data[13]), .B(idata[13]), .S0(n694), .Y(n481) );
  MX2XL U607 ( .A(data[14]), .B(idata[14]), .S0(n694), .Y(n482) );
  MX2XL U608 ( .A(data[15]), .B(idata[15]), .S0(n694), .Y(n483) );
  MX2XL U609 ( .A(data[16]), .B(idata[16]), .S0(n694), .Y(n484) );
  MX2XL U610 ( .A(data[17]), .B(idata[17]), .S0(n694), .Y(n485) );
  MX2XL U611 ( .A(data[18]), .B(idata[18]), .S0(n694), .Y(n486) );
  CLKBUFX3 U612 ( .A(n1125), .Y(n679) );
  CLKBUFX3 U613 ( .A(n1124), .Y(n677) );
  CLKBUFX3 U614 ( .A(n1121), .Y(n671) );
  CLKBUFX3 U615 ( .A(n1123), .Y(n675) );
  CLKBUFX3 U616 ( .A(n1122), .Y(n673) );
  AND2X2 U617 ( .A(n595), .B(n596), .Y(n594) );
  CLKINVX1 U618 ( .A(n742), .Y(n738) );
  OAI31X1 U619 ( .A0(n781), .A1(n812), .A2(n779), .B0(n695), .Y(n739) );
  NAND2X1 U620 ( .A(n816), .B(n695), .Y(n733) );
  NAND2X1 U621 ( .A(n695), .B(n779), .Y(n737) );
  NAND2X1 U622 ( .A(n695), .B(n781), .Y(n732) );
  NAND2X1 U623 ( .A(n695), .B(n780), .Y(n742) );
  NAND2X1 U624 ( .A(n598), .B(n721), .Y(n724) );
  CLKINVX1 U625 ( .A(n816), .Y(n721) );
  AOI21X1 U626 ( .A0(n695), .A1(n782), .B0(n738), .Y(n595) );
  AOI21X1 U627 ( .A0(n695), .A1(n726), .B0(n597), .Y(n596) );
  CLKBUFX3 U628 ( .A(n740), .Y(n693) );
  NOR2BX1 U629 ( .AN(n695), .B(n814), .Y(n597) );
  CLKBUFX3 U630 ( .A(n740), .Y(n695) );
  CLKBUFX3 U631 ( .A(n774), .Y(n699) );
  CLKBUFX3 U632 ( .A(n774), .Y(n698) );
  CLKBUFX3 U633 ( .A(n716), .Y(n707) );
  CLKBUFX3 U634 ( .A(n701), .Y(n706) );
  CLKBUFX3 U635 ( .A(n700), .Y(n713) );
  CLKBUFX3 U636 ( .A(n702), .Y(n714) );
  CLKBUFX3 U637 ( .A(n715), .Y(n711) );
  CLKBUFX3 U638 ( .A(n700), .Y(n712) );
  CLKBUFX3 U639 ( .A(n717), .Y(n705) );
  CLKBUFX3 U640 ( .A(n716), .Y(n708) );
  CLKBUFX3 U641 ( .A(n716), .Y(n709) );
  CLKBUFX3 U642 ( .A(n715), .Y(n710) );
  CLKBUFX3 U643 ( .A(n717), .Y(n704) );
  NAND2X1 U644 ( .A(n695), .B(n725), .Y(n735) );
  CLKINVX1 U645 ( .A(n813), .Y(n725) );
  NOR2X4 U646 ( .A(n665), .B(n898), .Y(n840) );
  CLKBUFX3 U647 ( .A(n841), .Y(n662) );
  NOR2X1 U648 ( .A(n811), .B(n665), .Y(n841) );
  CLKINVX1 U649 ( .A(n895), .Y(n779) );
  CLKINVX1 U650 ( .A(n898), .Y(n781) );
  CLKBUFX3 U651 ( .A(n845), .Y(n658) );
  NOR2X1 U652 ( .A(n894), .B(n665), .Y(n845) );
  CLKINVX1 U653 ( .A(n810), .Y(n782) );
  CLKBUFX3 U654 ( .A(n843), .Y(n663) );
  NOR2X1 U655 ( .A(n665), .B(n810), .Y(n843) );
  CLKBUFX3 U656 ( .A(n846), .Y(n657) );
  NOR2X1 U657 ( .A(n665), .B(n815), .Y(n846) );
  CLKINVX1 U658 ( .A(n896), .Y(n812) );
  AND2X2 U659 ( .A(n896), .B(n811), .Y(n598) );
  CLKBUFX3 U660 ( .A(n773), .Y(n697) );
  CLKBUFX3 U661 ( .A(n773), .Y(n696) );
  CLKBUFX3 U662 ( .A(n842), .Y(n664) );
  NOR2X1 U663 ( .A(n665), .B(n813), .Y(n842) );
  CLKBUFX3 U664 ( .A(n844), .Y(n659) );
  NOR2X1 U665 ( .A(n665), .B(n895), .Y(n844) );
  CLKINVX1 U666 ( .A(n897), .Y(n780) );
  CLKINVX1 U667 ( .A(n815), .Y(n726) );
  AO21X1 U668 ( .A0(n815), .A1(n896), .B0(n731), .Y(n734) );
  CLKBUFX3 U669 ( .A(n847), .Y(n661) );
  NOR2X1 U670 ( .A(n665), .B(n897), .Y(n847) );
  CLKBUFX3 U671 ( .A(n848), .Y(n660) );
  NOR2X1 U672 ( .A(n896), .B(n665), .Y(n848) );
  INVX3 U673 ( .A(n665), .Y(n853) );
  CLKINVX1 U674 ( .A(\sub_62/carry[10] ), .Y(n645) );
  CLKINVX1 U675 ( .A(n756), .Y(n751) );
  CLKINVX1 U676 ( .A(n765), .Y(n762) );
  CLKBUFX3 U677 ( .A(n701), .Y(n716) );
  CLKBUFX3 U678 ( .A(n700), .Y(n715) );
  CLKBUFX3 U679 ( .A(n701), .Y(n717) );
  NAND3BX1 U680 ( .AN(n746), .B(n947), .C(n667), .Y(n754) );
  NAND3BX1 U681 ( .AN(n946), .B(n667), .C(n746), .Y(n753) );
  AND2X2 U682 ( .A(n667), .B(n948), .Y(n907) );
  XNOR2X1 U683 ( .A(n673), .B(\sub_62/carry[9] ), .Y(N172) );
  XNOR2X1 U684 ( .A(n671), .B(\sub_62/carry[10] ), .Y(N173) );
  XNOR2X1 U685 ( .A(n692), .B(\sub_62/carry[11] ), .Y(N174) );
  NAND2X1 U686 ( .A(n647), .B(n645), .Y(\sub_62/carry[11] ) );
  XNOR2X1 U687 ( .A(n683), .B(\sub_54/carry[4] ), .Y(N142) );
  XNOR2X1 U688 ( .A(n681), .B(\sub_54/carry[5] ), .Y(N143) );
  XOR2X1 U689 ( .A(n679), .B(\sub_54/carry[6] ), .Y(N144) );
  XOR2X1 U690 ( .A(n677), .B(n679), .Y(N424) );
  XNOR2X1 U691 ( .A(n677), .B(n679), .Y(N157) );
  XNOR2X1 U692 ( .A(n677), .B(n603), .Y(N145) );
  XNOR2X1 U693 ( .A(n689), .B(caddr_wr[0]), .Y(N139) );
  XNOR2X1 U694 ( .A(n687), .B(\sub_54/carry[2] ), .Y(N140) );
  XNOR2X1 U695 ( .A(n685), .B(\sub_54/carry[3] ), .Y(N141) );
  OAI31X1 U696 ( .A0(n724), .A1(n780), .A2(n726), .B0(n1106), .Y(n731) );
  XNOR2X1 U697 ( .A(n675), .B(\sub_62/carry[8] ), .Y(N171) );
  OAI211X1 U698 ( .A0(n898), .A1(n960), .B0(n831), .C0(n810), .Y(n720) );
  AOI31X1 U699 ( .A0(n814), .A1(n957), .A2(n958), .B0(n802), .Y(n719) );
  OAI22XL U700 ( .A0(n895), .A1(n778), .B0(n963), .B1(n964), .Y(n718) );
  OAI31XL U701 ( .A0(n724), .A1(n780), .A2(n538), .B0(n699), .Y(n722) );
  CLKINVX1 U702 ( .A(n961), .Y(n778) );
  OAI21XL U703 ( .A0(n899), .A1(n900), .B0(n1106), .Y(n837) );
  CLKINVX1 U704 ( .A(caddr_wr[0]), .Y(N470) );
  CLKINVX1 U705 ( .A(n811), .Y(n954) );
  CLKBUFX3 U706 ( .A(n818), .Y(n655) );
  OAI21XL U707 ( .A0(n830), .A1(n801), .B0(n656), .Y(n818) );
  NAND2X1 U708 ( .A(n752), .B(n1077), .Y(n756) );
  NAND2X1 U709 ( .A(n759), .B(n1082), .Y(n764) );
  NAND2X1 U710 ( .A(n760), .B(n1082), .Y(n765) );
  AND2X2 U711 ( .A(n668), .B(n808), .Y(n971) );
  AND2X2 U712 ( .A(n668), .B(n996), .Y(n972) );
  AND3X2 U713 ( .A(n668), .B(n997), .C(n1000), .Y(n973) );
  XNOR2X1 U714 ( .A(n692), .B(\sub_54/carry[11] ), .Y(N149) );
  NAND2X1 U715 ( .A(n647), .B(n648), .Y(\sub_54/carry[11] ) );
  CLKINVX1 U716 ( .A(n671), .Y(n647) );
  CLKINVX1 U717 ( .A(\sub_54/carry[10] ), .Y(n648) );
  OR2X1 U718 ( .A(n689), .B(caddr_wr[0]), .Y(\sub_54/carry[2] ) );
  OR2X1 U719 ( .A(n687), .B(\sub_54/carry[2] ), .Y(\sub_54/carry[3] ) );
  OR2X1 U720 ( .A(n677), .B(n603), .Y(\sub_54/carry[8] ) );
  OR2X1 U721 ( .A(n675), .B(\sub_54/carry[8] ), .Y(\sub_54/carry[9] ) );
  OR2X1 U722 ( .A(n683), .B(\sub_54/carry[4] ), .Y(\sub_54/carry[5] ) );
  OR2X1 U723 ( .A(n673), .B(\sub_54/carry[9] ), .Y(\sub_54/carry[10] ) );
  OR2X1 U724 ( .A(n681), .B(\sub_54/carry[5] ), .Y(\sub_54/carry[6] ) );
  AND2X2 U725 ( .A(n642), .B(n769), .Y(n599) );
  AND2X2 U726 ( .A(n601), .B(n641), .Y(n600) );
  AND2X2 U727 ( .A(n642), .B(n767), .Y(n601) );
  AND2X2 U728 ( .A(n640), .B(n756), .Y(n602) );
  AND2X2 U729 ( .A(n679), .B(\sub_54/carry[6] ), .Y(n603) );
  AND2X2 U730 ( .A(n641), .B(n599), .Y(n604) );
  CLKINVX1 U731 ( .A(n761), .Y(n759) );
  CLKINVX1 U732 ( .A(n763), .Y(n760) );
  OR2X1 U733 ( .A(n685), .B(\sub_54/carry[3] ), .Y(\sub_54/carry[4] ) );
  XNOR2X1 U734 ( .A(n677), .B(\sub_62/carry[7] ), .Y(N170) );
  XOR2X1 U735 ( .A(n677), .B(\add_103/carry[7] ), .Y(N477) );
  XNOR2X1 U736 ( .A(n675), .B(\sub_54/carry[8] ), .Y(N146) );
  XNOR2X1 U737 ( .A(n673), .B(\sub_54/carry[9] ), .Y(N147) );
  XNOR2X1 U738 ( .A(n671), .B(\sub_54/carry[10] ), .Y(N148) );
  XOR2X1 U739 ( .A(n679), .B(\add_90/carry[6] ), .Y(N370) );
  XOR2X1 U740 ( .A(n675), .B(n608), .Y(N478) );
  XOR2X1 U741 ( .A(n673), .B(n620), .Y(N479) );
  XOR2X1 U742 ( .A(n671), .B(n621), .Y(N480) );
  XNOR2X1 U743 ( .A(n692), .B(n650), .Y(N481) );
  NAND2X1 U744 ( .A(n671), .B(n621), .Y(n650) );
  XOR2X1 U745 ( .A(n677), .B(n607), .Y(N371) );
  XOR2X1 U746 ( .A(n675), .B(n611), .Y(N372) );
  XOR2X1 U747 ( .A(n673), .B(n612), .Y(N373) );
  XOR2X1 U748 ( .A(n671), .B(n613), .Y(N374) );
  CLKINVX1 U749 ( .A(n965), .Y(n960) );
  OR2X1 U750 ( .A(n689), .B(caddr_wr[0]), .Y(\add_90/carry[2] ) );
  OR2X1 U751 ( .A(n687), .B(\add_90/carry[2] ), .Y(\add_90/carry[3] ) );
  OR2X1 U752 ( .A(n685), .B(\add_90/carry[3] ), .Y(\add_90/carry[4] ) );
  OR2X1 U753 ( .A(n683), .B(\add_90/carry[4] ), .Y(\add_90/carry[5] ) );
  OR2X1 U754 ( .A(n679), .B(n609), .Y(\sub_62/carry[7] ) );
  OR2X1 U755 ( .A(n677), .B(\sub_62/carry[7] ), .Y(\sub_62/carry[8] ) );
  OR2X1 U756 ( .A(n675), .B(\sub_62/carry[8] ), .Y(\sub_62/carry[9] ) );
  OR2X1 U757 ( .A(n673), .B(\sub_62/carry[9] ), .Y(\sub_62/carry[10] ) );
  OR2X1 U758 ( .A(n681), .B(\add_90/carry[5] ), .Y(\add_90/carry[6] ) );
  OR2X1 U759 ( .A(n679), .B(n610), .Y(\add_103/carry[7] ) );
  AND2X2 U760 ( .A(n689), .B(caddr_wr[0]), .Y(n605) );
  AND2X2 U761 ( .A(n689), .B(caddr_wr[0]), .Y(n606) );
  AND2X2 U762 ( .A(n679), .B(\add_90/carry[6] ), .Y(n607) );
  AND2X2 U763 ( .A(n677), .B(\add_103/carry[7] ), .Y(n608) );
  AND2X2 U764 ( .A(n681), .B(n618), .Y(n609) );
  AND2X2 U765 ( .A(n681), .B(n619), .Y(n610) );
  AND2X2 U766 ( .A(n677), .B(n607), .Y(n611) );
  AND2X2 U767 ( .A(n675), .B(n611), .Y(n612) );
  AND2X2 U768 ( .A(n673), .B(n612), .Y(n613) );
  AND2X2 U769 ( .A(n687), .B(n605), .Y(n614) );
  AND2X2 U770 ( .A(n687), .B(n606), .Y(n615) );
  AND2X2 U771 ( .A(n685), .B(n614), .Y(n616) );
  AND2X2 U772 ( .A(n685), .B(n615), .Y(n617) );
  AND2X2 U773 ( .A(n683), .B(n616), .Y(n618) );
  AND2X2 U774 ( .A(n683), .B(n617), .Y(n619) );
  AND2X2 U775 ( .A(n675), .B(n608), .Y(n620) );
  AND2X2 U776 ( .A(n673), .B(n620), .Y(n621) );
  OAI2BB1X1 U777 ( .A0N(n644), .A1N(n636), .B0(n767), .Y(N620) );
  CLKINVX1 U778 ( .A(n769), .Y(n766) );
  XNOR2X1 U779 ( .A(n692), .B(n652), .Y(N375) );
  NAND2X1 U780 ( .A(n671), .B(n613), .Y(n652) );
  XNOR2X1 U781 ( .A(n689), .B(caddr_wr[0]), .Y(N365) );
  XNOR2X1 U782 ( .A(n679), .B(n609), .Y(N169) );
  XNOR2X1 U783 ( .A(n687), .B(\add_90/carry[2] ), .Y(N366) );
  XNOR2X1 U784 ( .A(n683), .B(\add_90/carry[4] ), .Y(N368) );
  XNOR2X1 U785 ( .A(n681), .B(\add_90/carry[5] ), .Y(N369) );
  XNOR2X1 U786 ( .A(n685), .B(\add_90/carry[3] ), .Y(N367) );
  XNOR2X1 U787 ( .A(n675), .B(\sub_57/carry[8] ), .Y(N158) );
  XNOR2X1 U788 ( .A(n673), .B(\sub_57/carry[9] ), .Y(N159) );
  XNOR2X1 U789 ( .A(n671), .B(\sub_57/carry[10] ), .Y(N160) );
  XNOR2X1 U790 ( .A(n679), .B(n610), .Y(N476) );
  XOR2X1 U791 ( .A(n687), .B(n605), .Y(N165) );
  XOR2X1 U792 ( .A(n683), .B(n616), .Y(N167) );
  XOR2X1 U793 ( .A(n681), .B(n618), .Y(N168) );
  XOR2X1 U794 ( .A(n685), .B(n614), .Y(N166) );
  XOR2X1 U795 ( .A(n687), .B(n606), .Y(N472) );
  XOR2X1 U796 ( .A(n683), .B(n617), .Y(N474) );
  XOR2X1 U797 ( .A(n681), .B(n619), .Y(N475) );
  XOR2X1 U798 ( .A(n685), .B(n615), .Y(N473) );
  XNOR2X1 U799 ( .A(n692), .B(\sub_57/carry[11] ), .Y(N161) );
  NAND2X1 U800 ( .A(n647), .B(n646), .Y(\sub_57/carry[11] ) );
  CLKINVX1 U801 ( .A(\sub_57/carry[10] ), .Y(n646) );
  XOR2X1 U802 ( .A(n675), .B(n622), .Y(N425) );
  XOR2X1 U803 ( .A(n673), .B(n623), .Y(N426) );
  XOR2X1 U804 ( .A(n671), .B(n624), .Y(N427) );
  XNOR2X1 U805 ( .A(n692), .B(n651), .Y(N428) );
  NAND2X1 U806 ( .A(n671), .B(n624), .Y(n651) );
  OR2X1 U807 ( .A(n677), .B(n679), .Y(\sub_57/carry[8] ) );
  OR2X1 U808 ( .A(n675), .B(\sub_57/carry[8] ), .Y(\sub_57/carry[9] ) );
  OR2X1 U809 ( .A(n673), .B(\sub_57/carry[9] ), .Y(\sub_57/carry[10] ) );
  AND2X2 U810 ( .A(n677), .B(n679), .Y(n622) );
  AND2X2 U811 ( .A(n675), .B(n622), .Y(n623) );
  AND2X2 U812 ( .A(n673), .B(n623), .Y(n624) );
  AO21X1 U813 ( .A0(n643), .A1(n602), .B0(n759), .Y(N616) );
  XOR2X1 U814 ( .A(n689), .B(caddr_wr[0]), .Y(N164) );
  XOR2X1 U815 ( .A(n689), .B(caddr_wr[0]), .Y(N471) );
  CLKBUFX3 U816 ( .A(n715), .Y(n703) );
  CLKBUFX3 U817 ( .A(n777), .Y(n702) );
  CLKBUFX3 U818 ( .A(n777), .Y(n700) );
  CLKBUFX3 U819 ( .A(n777), .Y(n701) );
  XOR2X1 U820 ( .A(N628), .B(N629), .Y(N609) );
  XOR2X1 U821 ( .A(n747), .B(N630), .Y(n748) );
  AOI2BB1X1 U822 ( .A0N(n1077), .A1N(n752), .B0(n751), .Y(n755) );
  XOR2X1 U823 ( .A(sum[20]), .B(sum[21]), .Y(N633) );
  XOR2X1 U824 ( .A(n1079), .B(n758), .Y(N634) );
  XOR2X1 U825 ( .A(sum[23]), .B(n638), .Y(N635) );
  AO21X1 U826 ( .A0(n643), .A1(n638), .B0(n760), .Y(N636) );
  AO21X1 U827 ( .A0(sum[25]), .A1(n763), .B0(n762), .Y(N637) );
  XOR2X1 U828 ( .A(n765), .B(sum[26]), .Y(N638) );
  XOR2X1 U829 ( .A(sum[27]), .B(n637), .Y(N639) );
  AO21X1 U830 ( .A0(n644), .A1(n637), .B0(n766), .Y(N640) );
  XOR2X1 U831 ( .A(n769), .B(sum[29]), .Y(N641) );
  XOR2X1 U832 ( .A(n1087), .B(n770), .Y(N642) );
  XOR2X1 U833 ( .A(sum[31]), .B(n599), .Y(N643) );
  XOR2X1 U834 ( .A(n1089), .B(n772), .Y(N644) );
  XOR2X1 U835 ( .A(sum[33]), .B(n604), .Y(N645) );
  XOR2X1 U836 ( .A(sum[34]), .B(n635), .Y(N646) );
  XOR2X1 U837 ( .A(n1092), .B(n745), .Y(N647) );
  BUFX16 U838 ( .A(N150), .Y(caddr_wr[0]) );
  OAI2BB2XL U839 ( .B0(n1093), .B1(n774), .A0N(N212), .A1N(n697), .Y(n464) );
  OAI2BB2XL U840 ( .B0(n1083), .B1(n698), .A0N(N202), .A1N(n697), .Y(n454) );
  OAI2BB2XL U841 ( .B0(n1086), .B1(n698), .A0N(N205), .A1N(n697), .Y(n457) );
  OAI2BB2XL U842 ( .B0(n1087), .B1(n698), .A0N(N206), .A1N(n697), .Y(n458) );
  OAI2BB2XL U843 ( .B0(n1095), .B1(n774), .A0N(N214), .A1N(n773), .Y(n466) );
  CLKBUFX3 U844 ( .A(N151), .Y(n689) );
  OAI2BB2XL U845 ( .B0(n1084), .B1(n698), .A0N(N203), .A1N(n697), .Y(n455) );
  XOR2XL U846 ( .A(n1149), .B(n629), .Y(N702) );
  XOR2XL U847 ( .A(n1150), .B(n628), .Y(N701) );
  XOR2XL U848 ( .A(n1148), .B(n630), .Y(N703) );
  XOR2X1 U849 ( .A(n1034), .B(n649), .Y(N704) );
  XNOR2XL U850 ( .A(n1149), .B(\sub_172/carry[9] ), .Y(N743) );
  XNOR2XL U851 ( .A(n1150), .B(\sub_172/carry[8] ), .Y(N742) );
  XNOR2XL U852 ( .A(n1148), .B(\sub_172/carry[10] ), .Y(N744) );
  XNOR2XL U853 ( .A(n1147), .B(\sub_172/carry[11] ), .Y(N745) );
  XOR2X1 U854 ( .A(n790), .B(n82), .Y(n535) );
  OAI211X1 U855 ( .A0(n1023), .A1(n694), .B0(n595), .C0(n735), .Y(n517) );
  OAI211X1 U856 ( .A0(n693), .A1(n541), .B0(n737), .C0(n594), .Y(n518) );
  OAI211X1 U857 ( .A0(n1029), .A1(n694), .B0(n733), .C0(n734), .Y(n527) );
  OAI211X1 U858 ( .A0(n1028), .A1(n695), .B0(n732), .C0(n735), .Y(n526) );
  OAI211X1 U859 ( .A0(n52), .A1(n694), .B0(n595), .C0(n739), .Y(n525) );
  OAI211X1 U860 ( .A0(n1027), .A1(n695), .B0(n734), .C0(n737), .Y(n524) );
  OAI211X1 U861 ( .A0(n1026), .A1(n694), .B0(n732), .C0(n742), .Y(n523) );
  NAND2X1 U862 ( .A(n739), .B(n730), .Y(n522) );
  CLKMX2X2 U863 ( .A(n539), .B(n810), .S0(n693), .Y(n730) );
  NAND4X1 U864 ( .A(n626), .B(n735), .C(n734), .D(n737), .Y(n529) );
  OAI2BB2XL U865 ( .B0(n1074), .B1(n698), .A0N(N193), .A1N(n696), .Y(n445) );
  OAI2BB2XL U866 ( .B0(n1080), .B1(n698), .A0N(N199), .A1N(n697), .Y(n451) );
  OAI2BB2XL U867 ( .B0(n1082), .B1(n698), .A0N(N201), .A1N(n697), .Y(n453) );
  NAND4X1 U868 ( .A(n595), .B(n732), .C(n737), .D(n729), .Y(n521) );
  AOI2BB1X1 U869 ( .A0N(n1025), .A1N(n695), .B0(n597), .Y(n729) );
  NAND3BX1 U870 ( .AN(n738), .B(n737), .C(n736), .Y(n530) );
  CLKMX2X2 U871 ( .A(n540), .B(n815), .S0(n693), .Y(n736) );
  OAI21XL U872 ( .A0(n1022), .A1(n693), .B0(n733), .Y(n515) );
  OAI21XL U873 ( .A0(n1021), .A1(n693), .B0(n733), .Y(n514) );
  OAI21XL U874 ( .A0(n1020), .A1(n693), .B0(n733), .Y(n513) );
  OAI21XL U875 ( .A0(n1019), .A1(n693), .B0(n733), .Y(n512) );
  NAND4BX1 U876 ( .AN(n727), .B(n735), .C(n596), .D(n739), .Y(n516) );
  NOR2X1 U877 ( .A(n693), .B(n51), .Y(n727) );
  AO22X1 U878 ( .A0(N191), .A1(n697), .B0(sum[15]), .B1(n723), .Y(n443) );
  NAND4X1 U879 ( .A(n728), .B(n735), .C(n594), .D(n732), .Y(n520) );
  MXI2X1 U880 ( .A(n1024), .B(n598), .S0(n693), .Y(n519) );
  NAND3X1 U881 ( .A(n739), .B(n742), .C(n741), .Y(n531) );
  OAI2BB2XL U882 ( .B0(n1039), .B1(n699), .A0N(N176), .A1N(n773), .Y(n408) );
  OAI2BB2XL U883 ( .B0(n1040), .B1(n699), .A0N(N177), .A1N(n773), .Y(n409) );
  OAI2BB2XL U884 ( .B0(n1041), .B1(n699), .A0N(N178), .A1N(n773), .Y(n410) );
  OAI2BB2XL U885 ( .B0(n1042), .B1(n699), .A0N(N179), .A1N(n696), .Y(n411) );
  OAI2BB2XL U886 ( .B0(n1043), .B1(n699), .A0N(N180), .A1N(n697), .Y(n412) );
  OAI2BB2XL U887 ( .B0(n1044), .B1(n699), .A0N(N181), .A1N(n696), .Y(n413) );
  OAI2BB2XL U888 ( .B0(n1045), .B1(n699), .A0N(N182), .A1N(n696), .Y(n414) );
  OAI2BB2XL U889 ( .B0(n1046), .B1(n698), .A0N(N183), .A1N(n696), .Y(n415) );
  OAI2BB2XL U890 ( .B0(n1047), .B1(n698), .A0N(N184), .A1N(n696), .Y(n416) );
  OAI2BB2XL U891 ( .B0(n1048), .B1(n698), .A0N(N185), .A1N(n696), .Y(n417) );
  OAI2BB2XL U892 ( .B0(n1049), .B1(n698), .A0N(N186), .A1N(n696), .Y(n418) );
  OAI2BB2XL U893 ( .B0(n1050), .B1(n698), .A0N(N187), .A1N(n696), .Y(n419) );
  OAI2BB2XL U894 ( .B0(n1051), .B1(n699), .A0N(N188), .A1N(n696), .Y(n420) );
  OAI2BB2XL U895 ( .B0(n1052), .B1(n698), .A0N(N189), .A1N(n696), .Y(n421) );
  OAI2BB2XL U896 ( .B0(n1053), .B1(n699), .A0N(N190), .A1N(n696), .Y(n422) );
  OAI2BB2XL U897 ( .B0(n1073), .B1(n698), .A0N(N192), .A1N(n696), .Y(n444) );
  OAI2BB2XL U898 ( .B0(n1075), .B1(n698), .A0N(N194), .A1N(n696), .Y(n446) );
  OAI2BB2XL U899 ( .B0(n1076), .B1(n774), .A0N(N195), .A1N(n696), .Y(n447) );
  OAI2BB2XL U900 ( .B0(n1077), .B1(n698), .A0N(N196), .A1N(n697), .Y(n448) );
  OAI2BB2XL U901 ( .B0(n1079), .B1(n698), .A0N(N198), .A1N(n697), .Y(n450) );
  OAI2BB2XL U902 ( .B0(n1081), .B1(n698), .A0N(N200), .A1N(n697), .Y(n452) );
  OAI21XL U903 ( .A0(n1030), .A1(n693), .B0(n596), .Y(n528) );
  CLKBUFX3 U904 ( .A(N152), .Y(n687) );
  CLKBUFX3 U905 ( .A(N153), .Y(n685) );
  CLKBUFX3 U906 ( .A(n817), .Y(n656) );
  AOI211X1 U907 ( .A0(n831), .A1(n832), .B0(n833), .C0(n82), .Y(n817) );
  OAI2BB2XL U908 ( .B0(n1078), .B1(n698), .A0N(N197), .A1N(n697), .Y(n449) );
  XNOR2XL U909 ( .A(n1153), .B(\add_153/carry[5] ), .Y(N698) );
  XNOR2XL U910 ( .A(n1154), .B(\add_153/carry[4] ), .Y(N697) );
  XNOR2XL U911 ( .A(n1155), .B(\add_153/carry[3] ), .Y(N696) );
  XOR2XL U912 ( .A(n1151), .B(n627), .Y(N700) );
  XOR2XL U913 ( .A(n1152), .B(\add_153/carry[6] ), .Y(N699) );
  XNOR2XL U914 ( .A(n1151), .B(\sub_172/carry[7] ), .Y(N741) );
  XNOR2XL U915 ( .A(n1152), .B(n625), .Y(N740) );
  XOR2XL U916 ( .A(n1153), .B(n631), .Y(N739) );
  XOR2XL U917 ( .A(n1154), .B(n632), .Y(N738) );
  XOR2XL U918 ( .A(n1155), .B(n633), .Y(N737) );
  XOR2XL U919 ( .A(n1156), .B(n634), .Y(N736) );
  XOR2XL U920 ( .A(n1157), .B(n1158), .Y(N735) );
  NAND2X1 U921 ( .A(N631), .B(n750), .Y(n752) );
  XOR2X1 U922 ( .A(n1089), .B(n771), .Y(N624) );
  NAND2X1 U923 ( .A(n601), .B(sum[31]), .Y(n771) );
  XOR2X1 U924 ( .A(n1092), .B(n744), .Y(N627) );
  NAND2X1 U925 ( .A(n639), .B(sum[34]), .Y(n744) );
  XOR2X1 U926 ( .A(sum[31]), .B(n601), .Y(N623) );
  XOR2X1 U927 ( .A(sum[34]), .B(n639), .Y(N626) );
  XOR2X1 U928 ( .A(sum[33]), .B(n600), .Y(N625) );
  AO21X1 U929 ( .A0(n636), .A1(sum[27]), .B0(sum[28]), .Y(n767) );
  AO21X1 U930 ( .A0(sum[27]), .A1(n637), .B0(sum[28]), .Y(n769) );
  AND2X2 U931 ( .A(sum[33]), .B(n604), .Y(n635) );
  NAND2X1 U932 ( .A(sum[34]), .B(n635), .Y(n745) );
  AO21X1 U933 ( .A0(n602), .A1(sum[23]), .B0(sum[24]), .Y(n761) );
  AO21X1 U934 ( .A0(sum[23]), .A1(n638), .B0(sum[24]), .Y(n763) );
  AND2X2 U935 ( .A(sum[26]), .B(n764), .Y(n636) );
  AND2X2 U936 ( .A(sum[26]), .B(n765), .Y(n637) );
  AND2X2 U937 ( .A(sum[20]), .B(n640), .Y(n638) );
  CLKBUFX3 U938 ( .A(N154), .Y(n683) );
  CLKBUFX3 U939 ( .A(N155), .Y(n681) );
  CLKINVX1 U940 ( .A(n743), .Y(n750) );
  NAND3BX1 U941 ( .AN(n1075), .B(N629), .C(N628), .Y(n743) );
  CLKBUFX3 U942 ( .A(n968), .Y(n668) );
  AOI2BB1X1 U943 ( .A0N(n1002), .A1N(n948), .B0(n82), .Y(n968) );
  AND2X2 U944 ( .A(n600), .B(sum[33]), .Y(n639) );
  AND2X2 U945 ( .A(sum[21]), .B(sum[22]), .Y(n640) );
  XNOR2XL U946 ( .A(n1157), .B(n1158), .Y(N694) );
  XNOR2XL U947 ( .A(n1156), .B(\add_153/carry[2] ), .Y(N695) );
  NAND2BX1 U948 ( .AN(state[0]), .B(n786), .Y(n784) );
  XOR2X1 U949 ( .A(n767), .B(sum[29]), .Y(N621) );
  XOR2X1 U950 ( .A(n764), .B(sum[26]), .Y(N618) );
  XOR2X1 U951 ( .A(n1087), .B(n768), .Y(N622) );
  NAND2X1 U952 ( .A(sum[29]), .B(n767), .Y(n768) );
  XOR2X1 U953 ( .A(sum[27]), .B(n636), .Y(N619) );
  NAND2X1 U954 ( .A(sum[29]), .B(n769), .Y(n770) );
  NAND2X1 U955 ( .A(n599), .B(sum[31]), .Y(n772) );
  OAI2BB1X1 U956 ( .A0N(sum[25]), .A1N(n761), .B0(n764), .Y(N617) );
  XOR2X1 U957 ( .A(n756), .B(sum[21]), .Y(N613) );
  XOR2X1 U958 ( .A(n1079), .B(n757), .Y(N614) );
  NAND2X1 U959 ( .A(sum[21]), .B(n756), .Y(n757) );
  XOR2X1 U960 ( .A(sum[23]), .B(n602), .Y(N615) );
  AND2X2 U961 ( .A(sum[31]), .B(sum[32]), .Y(n641) );
  AND2X2 U962 ( .A(sum[29]), .B(sum[30]), .Y(n642) );
  CLKBUFX3 U963 ( .A(n1120), .Y(n692) );
  BUFX12 U964 ( .A(N151), .Y(caddr_wr[1]) );
  BUFX12 U965 ( .A(N152), .Y(caddr_wr[2]) );
  BUFX12 U966 ( .A(N153), .Y(caddr_wr[3]) );
  BUFX12 U967 ( .A(N154), .Y(caddr_wr[4]) );
  BUFX12 U968 ( .A(N155), .Y(caddr_wr[5]) );
  BUFX12 U969 ( .A(n1125), .Y(caddr_wr[6]) );
  BUFX12 U970 ( .A(n1124), .Y(caddr_wr[7]) );
  BUFX12 U971 ( .A(n1123), .Y(caddr_wr[8]) );
  BUFX12 U972 ( .A(n1122), .Y(caddr_wr[9]) );
  BUFX12 U973 ( .A(n1121), .Y(caddr_wr[10]) );
  BUFX12 U974 ( .A(n1120), .Y(caddr_wr[11]) );
  BUFX12 U975 ( .A(n1106), .Y(busy) );
  NAND2X1 U976 ( .A(sum[20]), .B(sum[21]), .Y(n758) );
  NAND2X1 U977 ( .A(N629), .B(N628), .Y(n747) );
  AND2X2 U978 ( .A(sum[24]), .B(sum[23]), .Y(n643) );
  AND2X2 U979 ( .A(sum[28]), .B(sum[27]), .Y(n644) );
  OA22XL U980 ( .A0(n754), .A1(n748), .B0(n1075), .B1(n753), .Y(n913) );
  OA22XL U981 ( .A0(n755), .A1(n754), .B0(sum[20]), .B1(n753), .Y(n917) );
  AOI21X4 U982 ( .A0(N705), .A1(n951), .B0(n952), .Y(n950) );
  AO21X4 U983 ( .A0(n654), .A1(N631), .B0(n653), .Y(n749) );
  OAI221X2 U984 ( .A0(n654), .A1(n752), .B0(N631), .B1(n750), .C0(n749), .Y(
        n915) );
  XOR2X1 U985 ( .A(\r406/carry[4] ), .B(state[4]), .Y(N940) );
  OAI211X1 U986 ( .A0(n783), .A1(n1106), .B0(n784), .C0(n785), .Y(n537) );
  OAI221XL U987 ( .A0(n785), .A1(n787), .B0(n788), .B1(n1106), .C0(n789), .Y(
        n536) );
  NAND2X1 U988 ( .A(N940), .B(n786), .Y(n789) );
  MXI2X1 U989 ( .A(n791), .B(ready), .S0(n82), .Y(n790) );
  OAI2BB1X1 U990 ( .A0N(N937), .A1N(n786), .B0(n792), .Y(n534) );
  MXI2X1 U991 ( .A(n793), .B(state[1]), .S0(n82), .Y(n792) );
  AO21X1 U992 ( .A0(N938), .A1(n786), .B0(n795), .Y(n533) );
  MXI2X1 U993 ( .A(n796), .B(n797), .S0(n82), .Y(n795) );
  AO21X1 U994 ( .A0(N939), .A1(n786), .B0(n798), .Y(n532) );
  MXI2X1 U995 ( .A(n796), .B(n799), .S0(n82), .Y(n798) );
  OA21XL U996 ( .A0(n800), .A1(n785), .B0(n794), .Y(n796) );
  NAND3X1 U997 ( .A(n801), .B(n778), .C(n802), .Y(n794) );
  AOI21X1 U998 ( .A0(n803), .A1(n804), .B0(n82), .Y(n786) );
  OAI21XL U999 ( .A0(n788), .A1(n799), .B0(n805), .Y(n804) );
  NAND2X1 U1000 ( .A(state[3]), .B(state[1]), .Y(n807) );
  OAI31XL U1001 ( .A0(n797), .A1(n808), .A2(n799), .B0(n788), .Y(n803) );
  NAND2X1 U1002 ( .A(n810), .B(n811), .Y(n809) );
  OAI22XL U1003 ( .A0(n55), .A1(n656), .B0(n655), .B1(n819), .Y(n511) );
  CLKINVX1 U1004 ( .A(N323), .Y(n819) );
  MXI2X1 U1005 ( .A(n656), .B(n655), .S0(n81), .Y(n510) );
  OAI22XL U1006 ( .A0(n80), .A1(n656), .B0(n655), .B1(n820), .Y(n509) );
  CLKINVX1 U1007 ( .A(N313), .Y(n820) );
  OAI22XL U1008 ( .A0(n79), .A1(n656), .B0(n655), .B1(n821), .Y(n508) );
  CLKINVX1 U1009 ( .A(N314), .Y(n821) );
  OAI22XL U1010 ( .A0(n78), .A1(n656), .B0(n655), .B1(n822), .Y(n507) );
  CLKINVX1 U1011 ( .A(N315), .Y(n822) );
  OAI22XL U1012 ( .A0(n77), .A1(n656), .B0(n655), .B1(n823), .Y(n506) );
  CLKINVX1 U1013 ( .A(N316), .Y(n823) );
  OAI22XL U1014 ( .A0(n76), .A1(n656), .B0(n655), .B1(n824), .Y(n505) );
  CLKINVX1 U1015 ( .A(N317), .Y(n824) );
  OAI22XL U1016 ( .A0(n72), .A1(n656), .B0(n655), .B1(n825), .Y(n504) );
  CLKINVX1 U1017 ( .A(N318), .Y(n825) );
  OAI22XL U1018 ( .A0(n71), .A1(n656), .B0(n655), .B1(n826), .Y(n503) );
  CLKINVX1 U1019 ( .A(N319), .Y(n826) );
  OAI22XL U1020 ( .A0(n70), .A1(n656), .B0(n655), .B1(n827), .Y(n502) );
  CLKINVX1 U1021 ( .A(N320), .Y(n827) );
  OAI22XL U1022 ( .A0(n69), .A1(n656), .B0(n655), .B1(n828), .Y(n501) );
  CLKINVX1 U1023 ( .A(N321), .Y(n828) );
  OAI22XL U1024 ( .A0(n68), .A1(n656), .B0(n655), .B1(n829), .Y(n500) );
  CLKINVX1 U1025 ( .A(N322), .Y(n829) );
  NAND3X1 U1026 ( .A(n834), .B(n835), .C(n836), .Y(n499) );
  CLKMX2X2 U1027 ( .A(n840), .B(n662), .S0(caddr_wr[0]), .Y(n839) );
  AO22X1 U1028 ( .A0(N470), .A1(n664), .B0(N470), .B1(n663), .Y(n838) );
  AOI222XL U1029 ( .A0(caddr_wr[0]), .A1(n659), .B0(N470), .B1(n658), .C0(
        caddr_wr[0]), .C1(n657), .Y(n835) );
  AOI22X1 U1030 ( .A0(N217), .A1(n661), .B0(N470), .B1(n660), .Y(n834) );
  NAND4X1 U1031 ( .A(n849), .B(n850), .C(n851), .D(n852), .Y(n498) );
  AOI222XL U1032 ( .A0(n689), .A1(n659), .B0(N139), .B1(n658), .C0(n689), .C1(
        n657), .Y(n852) );
  AOI22X1 U1033 ( .A0(N218), .A1(n661), .B0(N164), .B1(n660), .Y(n851) );
  AOI222XL U1034 ( .A0(N365), .A1(n663), .B0(n662), .B1(caddr_wr[1]), .C0(n840), .C1(N313), .Y(n850) );
  AOI2BB2X1 U1035 ( .B0(N471), .B1(n664), .A0N(n1018), .A1N(n853), .Y(n849) );
  NAND4X1 U1036 ( .A(n854), .B(n855), .C(n856), .D(n857), .Y(n497) );
  AOI222XL U1037 ( .A0(n687), .A1(n659), .B0(N140), .B1(n658), .C0(n687), .C1(
        n657), .Y(n857) );
  AOI22X1 U1038 ( .A0(N219), .A1(n661), .B0(N165), .B1(n660), .Y(n856) );
  AOI222XL U1039 ( .A0(N366), .A1(n663), .B0(n662), .B1(caddr_wr[2]), .C0(n840), .C1(N314), .Y(n855) );
  AOI2BB2X1 U1040 ( .B0(N472), .B1(n664), .A0N(n1017), .A1N(n853), .Y(n854) );
  NAND4X1 U1041 ( .A(n858), .B(n859), .C(n860), .D(n861), .Y(n496) );
  AOI222XL U1042 ( .A0(n685), .A1(n659), .B0(N141), .B1(n658), .C0(n685), .C1(
        n657), .Y(n861) );
  AOI22X1 U1043 ( .A0(N220), .A1(n661), .B0(N166), .B1(n660), .Y(n860) );
  AOI222XL U1044 ( .A0(N367), .A1(n663), .B0(n662), .B1(caddr_wr[3]), .C0(n840), .C1(N315), .Y(n859) );
  AOI2BB2X1 U1045 ( .B0(N473), .B1(n664), .A0N(n1016), .A1N(n853), .Y(n858) );
  NAND4X1 U1046 ( .A(n862), .B(n863), .C(n864), .D(n865), .Y(n495) );
  AOI222XL U1047 ( .A0(n683), .A1(n659), .B0(N142), .B1(n658), .C0(n683), .C1(
        n657), .Y(n865) );
  AOI22X1 U1048 ( .A0(N221), .A1(n661), .B0(N167), .B1(n660), .Y(n864) );
  AOI222XL U1049 ( .A0(N368), .A1(n663), .B0(n662), .B1(caddr_wr[4]), .C0(n840), .C1(N316), .Y(n863) );
  AOI2BB2X1 U1050 ( .B0(N474), .B1(n664), .A0N(n1104), .A1N(n853), .Y(n862) );
  NAND4X1 U1051 ( .A(n866), .B(n867), .C(n868), .D(n869), .Y(n494) );
  AOI222XL U1052 ( .A0(n681), .A1(n659), .B0(N143), .B1(n658), .C0(n681), .C1(
        n657), .Y(n869) );
  AOI22X1 U1053 ( .A0(N222), .A1(n661), .B0(N168), .B1(n660), .Y(n868) );
  AOI222XL U1054 ( .A0(N369), .A1(n663), .B0(n662), .B1(caddr_wr[5]), .C0(n840), .C1(N317), .Y(n867) );
  AOI2BB2X1 U1055 ( .B0(N475), .B1(n664), .A0N(n1103), .A1N(n853), .Y(n866) );
  NAND4X1 U1056 ( .A(n870), .B(n871), .C(n872), .D(n873), .Y(n493) );
  AOI222XL U1057 ( .A0(n72), .A1(n659), .B0(N144), .B1(n658), .C0(n72), .C1(
        n657), .Y(n873) );
  AOI22X1 U1058 ( .A0(N223), .A1(n661), .B0(N169), .B1(n660), .Y(n872) );
  AOI222XL U1059 ( .A0(N370), .A1(n663), .B0(n662), .B1(caddr_wr[6]), .C0(n840), .C1(N318), .Y(n871) );
  AOI2BB2X1 U1060 ( .B0(N476), .B1(n664), .A0N(n1102), .A1N(n853), .Y(n870) );
  NAND4X1 U1061 ( .A(n874), .B(n875), .C(n876), .D(n877), .Y(n492) );
  AOI222XL U1062 ( .A0(N424), .A1(n659), .B0(N145), .B1(n658), .C0(N157), .C1(
        n657), .Y(n877) );
  AOI22X1 U1063 ( .A0(N224), .A1(n661), .B0(N170), .B1(n660), .Y(n876) );
  AOI222XL U1064 ( .A0(N371), .A1(n663), .B0(n662), .B1(caddr_wr[7]), .C0(n840), .C1(N319), .Y(n875) );
  AOI2BB2X1 U1065 ( .B0(N477), .B1(n664), .A0N(n1101), .A1N(n853), .Y(n874) );
  NAND4X1 U1066 ( .A(n878), .B(n879), .C(n880), .D(n881), .Y(n491) );
  AOI222XL U1067 ( .A0(N425), .A1(n659), .B0(N146), .B1(n658), .C0(N158), .C1(
        n657), .Y(n881) );
  AOI22X1 U1068 ( .A0(N225), .A1(n661), .B0(N171), .B1(n660), .Y(n880) );
  AOI222XL U1069 ( .A0(N372), .A1(n663), .B0(n662), .B1(caddr_wr[8]), .C0(n840), .C1(N320), .Y(n879) );
  AOI2BB2X1 U1070 ( .B0(N478), .B1(n664), .A0N(n1100), .A1N(n853), .Y(n878) );
  NAND4X1 U1071 ( .A(n882), .B(n883), .C(n884), .D(n885), .Y(n490) );
  AOI222XL U1072 ( .A0(N426), .A1(n659), .B0(N147), .B1(n658), .C0(N159), .C1(
        n657), .Y(n885) );
  AOI22X1 U1073 ( .A0(N226), .A1(n661), .B0(N172), .B1(n660), .Y(n884) );
  AOI222XL U1074 ( .A0(N373), .A1(n663), .B0(n662), .B1(caddr_wr[9]), .C0(n840), .C1(N321), .Y(n883) );
  AOI2BB2X1 U1075 ( .B0(N479), .B1(n664), .A0N(n1099), .A1N(n853), .Y(n882) );
  NAND4X1 U1076 ( .A(n886), .B(n887), .C(n888), .D(n889), .Y(n489) );
  AOI222XL U1077 ( .A0(N427), .A1(n659), .B0(N148), .B1(n658), .C0(N160), .C1(
        n657), .Y(n889) );
  AOI22X1 U1078 ( .A0(N227), .A1(n661), .B0(N173), .B1(n660), .Y(n888) );
  AOI222XL U1079 ( .A0(N374), .A1(n663), .B0(n662), .B1(caddr_wr[10]), .C0(
        n840), .C1(N322), .Y(n887) );
  AOI2BB2X1 U1080 ( .B0(N480), .B1(n664), .A0N(n1098), .A1N(n853), .Y(n886) );
  NAND4X1 U1081 ( .A(n890), .B(n891), .C(n892), .D(n893), .Y(n488) );
  AOI222XL U1082 ( .A0(N428), .A1(n659), .B0(N149), .B1(n658), .C0(N161), .C1(
        n657), .Y(n893) );
  AOI22X1 U1083 ( .A0(N228), .A1(n661), .B0(N174), .B1(n660), .Y(n892) );
  AOI222XL U1084 ( .A0(N375), .A1(n663), .B0(n662), .B1(caddr_wr[11]), .C0(
        n840), .C1(N323), .Y(n891) );
  AOI2BB2X1 U1085 ( .B0(N481), .B1(n664), .A0N(n1097), .A1N(n853), .Y(n890) );
  NAND3X1 U1086 ( .A(n901), .B(n894), .C(n598), .Y(n900) );
  NAND3X1 U1087 ( .A(n897), .B(n815), .C(n813), .Y(n899) );
  NAND2X1 U1088 ( .A(n902), .B(n903), .Y(n815) );
  OAI211X1 U1089 ( .A0(n104), .A1(n667), .B0(n905), .C0(n906), .Y(n442) );
  AOI22X1 U1090 ( .A0(N627), .A1(n653), .B0(N647), .B1(n654), .Y(n906) );
  NAND2X1 U1091 ( .A(cdata_rd[19]), .B(n666), .Y(n905) );
  OAI211X1 U1092 ( .A0(n1072), .A1(n667), .B0(n908), .C0(n909), .Y(n441) );
  AOI22X1 U1093 ( .A0(n1073), .A1(n653), .B0(N628), .B1(n654), .Y(n909) );
  NAND2X1 U1094 ( .A(cdata_rd[0]), .B(n666), .Y(n908) );
  OAI211X1 U1095 ( .A0(n1071), .A1(n667), .B0(n910), .C0(n911), .Y(n440) );
  AOI22X1 U1096 ( .A0(N609), .A1(n653), .B0(N629), .B1(n654), .Y(n911) );
  NAND2X1 U1097 ( .A(cdata_rd[1]), .B(n666), .Y(n910) );
  OAI211X1 U1098 ( .A0(n1070), .A1(n667), .B0(n912), .C0(n913), .Y(n439) );
  OAI211X1 U1099 ( .A0(n1069), .A1(n667), .B0(n914), .C0(n915), .Y(n438) );
  NAND2X1 U1100 ( .A(cdata_rd[3]), .B(n666), .Y(n914) );
  OAI211X1 U1101 ( .A0(n1068), .A1(n667), .B0(n916), .C0(n917), .Y(n437) );
  NAND2X1 U1102 ( .A(cdata_rd[4]), .B(n666), .Y(n916) );
  OAI211X1 U1103 ( .A0(n1067), .A1(n667), .B0(n918), .C0(n919), .Y(n436) );
  AOI22X1 U1104 ( .A0(N613), .A1(n653), .B0(N633), .B1(n654), .Y(n919) );
  NAND2X1 U1105 ( .A(cdata_rd[5]), .B(n666), .Y(n918) );
  OAI211X1 U1106 ( .A0(n1066), .A1(n667), .B0(n920), .C0(n921), .Y(n435) );
  AOI22X1 U1107 ( .A0(N614), .A1(n653), .B0(N634), .B1(n654), .Y(n921) );
  NAND2X1 U1108 ( .A(cdata_rd[6]), .B(n666), .Y(n920) );
  OAI211X1 U1109 ( .A0(n1065), .A1(n667), .B0(n922), .C0(n923), .Y(n434) );
  AOI22X1 U1110 ( .A0(N615), .A1(n653), .B0(N635), .B1(n654), .Y(n923) );
  NAND2X1 U1111 ( .A(cdata_rd[7]), .B(n666), .Y(n922) );
  OAI211X1 U1112 ( .A0(n1064), .A1(n667), .B0(n924), .C0(n925), .Y(n433) );
  AOI22X1 U1113 ( .A0(N616), .A1(n653), .B0(N636), .B1(n654), .Y(n925) );
  NAND2X1 U1114 ( .A(cdata_rd[8]), .B(n666), .Y(n924) );
  OAI211X1 U1115 ( .A0(n1063), .A1(n667), .B0(n926), .C0(n927), .Y(n432) );
  AOI22X1 U1116 ( .A0(N617), .A1(n653), .B0(N637), .B1(n654), .Y(n927) );
  NAND2X1 U1117 ( .A(cdata_rd[9]), .B(n666), .Y(n926) );
  OAI211X1 U1118 ( .A0(n1062), .A1(n667), .B0(n928), .C0(n929), .Y(n431) );
  AOI22X1 U1119 ( .A0(N618), .A1(n653), .B0(N638), .B1(n654), .Y(n929) );
  NAND2X1 U1120 ( .A(cdata_rd[10]), .B(n666), .Y(n928) );
  OAI211X1 U1121 ( .A0(n1061), .A1(n667), .B0(n930), .C0(n931), .Y(n430) );
  AOI22X1 U1122 ( .A0(N619), .A1(n653), .B0(N639), .B1(n654), .Y(n931) );
  NAND2X1 U1123 ( .A(cdata_rd[11]), .B(n666), .Y(n930) );
  OAI211X1 U1124 ( .A0(n1060), .A1(n667), .B0(n932), .C0(n933), .Y(n429) );
  AOI22X1 U1125 ( .A0(N620), .A1(n653), .B0(N640), .B1(n654), .Y(n933) );
  NAND2X1 U1126 ( .A(cdata_rd[12]), .B(n666), .Y(n932) );
  OAI211X1 U1127 ( .A0(n1059), .A1(n667), .B0(n934), .C0(n935), .Y(n428) );
  AOI22X1 U1128 ( .A0(N621), .A1(n653), .B0(N641), .B1(n654), .Y(n935) );
  NAND2X1 U1129 ( .A(cdata_rd[13]), .B(n666), .Y(n934) );
  OAI211X1 U1130 ( .A0(n1058), .A1(n667), .B0(n936), .C0(n937), .Y(n427) );
  AOI22X1 U1131 ( .A0(N622), .A1(n653), .B0(N642), .B1(n654), .Y(n937) );
  NAND2X1 U1132 ( .A(cdata_rd[14]), .B(n666), .Y(n936) );
  OAI211X1 U1133 ( .A0(n1057), .A1(n667), .B0(n938), .C0(n939), .Y(n426) );
  AOI22X1 U1134 ( .A0(N623), .A1(n653), .B0(N643), .B1(n654), .Y(n939) );
  NAND2X1 U1135 ( .A(cdata_rd[15]), .B(n666), .Y(n938) );
  OAI211X1 U1136 ( .A0(n1056), .A1(n667), .B0(n940), .C0(n941), .Y(n425) );
  AOI22X1 U1137 ( .A0(N624), .A1(n653), .B0(N644), .B1(n654), .Y(n941) );
  NAND2X1 U1138 ( .A(cdata_rd[16]), .B(n666), .Y(n940) );
  OAI211X1 U1139 ( .A0(n1055), .A1(n667), .B0(n942), .C0(n943), .Y(n424) );
  AOI22X1 U1140 ( .A0(N625), .A1(n653), .B0(N645), .B1(n654), .Y(n943) );
  NAND2X1 U1141 ( .A(cdata_rd[17]), .B(n666), .Y(n942) );
  OAI211X1 U1142 ( .A0(n1054), .A1(n667), .B0(n944), .C0(n945), .Y(n423) );
  AOI22X1 U1143 ( .A0(N626), .A1(n653), .B0(N646), .B1(n654), .Y(n945) );
  NAND2X1 U1144 ( .A(cdata_rd[18]), .B(n666), .Y(n944) );
  NOR2BX1 U1145 ( .AN(n953), .B(n947), .Y(n949) );
  CLKINVX1 U1146 ( .A(n946), .Y(n947) );
  NAND3X1 U1147 ( .A(n814), .B(n813), .C(n901), .Y(n816) );
  NOR3X1 U1148 ( .A(n781), .B(n782), .C(n779), .Y(n901) );
  NAND2X1 U1149 ( .A(n955), .B(n956), .Y(n810) );
  NOR3BXL U1150 ( .AN(n959), .B(n55), .C(n68), .Y(n802) );
  OR2X1 U1151 ( .A(n813), .B(n960), .Y(n958) );
  NAND2X1 U1152 ( .A(n808), .B(n538), .Y(n813) );
  NAND2X1 U1153 ( .A(n538), .B(n903), .Y(n814) );
  NAND3X1 U1154 ( .A(n538), .B(n961), .C(n955), .Y(n957) );
  NAND2X1 U1155 ( .A(n956), .B(n903), .Y(n898) );
  NOR4X1 U1156 ( .A(n966), .B(n1125), .C(n1123), .D(n1124), .Y(n964) );
  NAND3X1 U1157 ( .A(n68), .B(n55), .C(n69), .Y(n966) );
  AOI221XL U1158 ( .A0(n812), .A1(n965), .B0(n954), .B1(n961), .C0(n780), .Y(
        n963) );
  NAND2X1 U1159 ( .A(n808), .B(n956), .Y(n811) );
  NAND4X1 U1160 ( .A(n79), .B(n78), .C(n80), .D(n967), .Y(n965) );
  NOR3X1 U1161 ( .A(N154), .B(N150), .C(N155), .Y(n967) );
  NAND2X1 U1162 ( .A(n902), .B(n955), .Y(n896) );
  NOR2BX1 U1163 ( .AN(n962), .B(state[3]), .Y(n902) );
  NOR2X1 U1164 ( .A(state[2]), .B(state[4]), .Y(n962) );
  NOR3X1 U1165 ( .A(state[3]), .B(state[4]), .C(n797), .Y(n956) );
  OAI211X1 U1166 ( .A0(n112), .A1(n668), .B0(n969), .C0(n970), .Y(n407) );
  AOI22X1 U1167 ( .A0(n112), .A1(n971), .B0(N681), .B1(n972), .Y(n970) );
  OAI211X1 U1168 ( .A0(n111), .A1(n668), .B0(n974), .C0(n975), .Y(n406) );
  AOI22X1 U1169 ( .A0(N694), .A1(n971), .B0(N682), .B1(n972), .Y(n975) );
  NAND2X1 U1170 ( .A(N735), .B(n973), .Y(n974) );
  OAI211X1 U1171 ( .A0(n110), .A1(n668), .B0(n976), .C0(n977), .Y(n405) );
  AOI22X1 U1172 ( .A0(N695), .A1(n971), .B0(N683), .B1(n972), .Y(n977) );
  NAND2X1 U1173 ( .A(N736), .B(n973), .Y(n976) );
  OAI211X1 U1174 ( .A0(n109), .A1(n668), .B0(n978), .C0(n979), .Y(n404) );
  AOI22X1 U1175 ( .A0(N696), .A1(n971), .B0(N684), .B1(n972), .Y(n979) );
  NAND2X1 U1176 ( .A(N737), .B(n973), .Y(n978) );
  OAI211X1 U1177 ( .A0(n108), .A1(n668), .B0(n980), .C0(n981), .Y(n403) );
  AOI22X1 U1178 ( .A0(N697), .A1(n971), .B0(N685), .B1(n972), .Y(n981) );
  NAND2X1 U1179 ( .A(N738), .B(n973), .Y(n980) );
  OAI211X1 U1180 ( .A0(n107), .A1(n668), .B0(n982), .C0(n983), .Y(n402) );
  AOI22X1 U1181 ( .A0(N698), .A1(n971), .B0(N686), .B1(n972), .Y(n983) );
  NAND2X1 U1182 ( .A(N739), .B(n973), .Y(n982) );
  OAI211X1 U1183 ( .A0(n106), .A1(n668), .B0(n984), .C0(n985), .Y(n401) );
  AOI22X1 U1184 ( .A0(N699), .A1(n971), .B0(N687), .B1(n972), .Y(n985) );
  NAND2X1 U1185 ( .A(N740), .B(n973), .Y(n984) );
  OAI211X1 U1186 ( .A0(n1038), .A1(n668), .B0(n986), .C0(n987), .Y(n400) );
  AOI22X1 U1187 ( .A0(N700), .A1(n971), .B0(N688), .B1(n972), .Y(n987) );
  NAND2X1 U1188 ( .A(N741), .B(n973), .Y(n986) );
  OAI211X1 U1189 ( .A0(n1037), .A1(n668), .B0(n988), .C0(n989), .Y(n399) );
  AOI22X1 U1190 ( .A0(N701), .A1(n971), .B0(N689), .B1(n972), .Y(n989) );
  NAND2X1 U1191 ( .A(N742), .B(n973), .Y(n988) );
  OAI211X1 U1192 ( .A0(n1036), .A1(n668), .B0(n990), .C0(n991), .Y(n398) );
  AOI22X1 U1193 ( .A0(N702), .A1(n971), .B0(N690), .B1(n972), .Y(n991) );
  NAND2X1 U1194 ( .A(N743), .B(n973), .Y(n990) );
  OAI211X1 U1195 ( .A0(n1035), .A1(n668), .B0(n992), .C0(n993), .Y(n397) );
  AOI22X1 U1196 ( .A0(N703), .A1(n971), .B0(N691), .B1(n972), .Y(n993) );
  NAND2X1 U1197 ( .A(N744), .B(n973), .Y(n992) );
  OAI211X1 U1198 ( .A0(n1034), .A1(n668), .B0(n994), .C0(n995), .Y(n396) );
  AOI22X1 U1199 ( .A0(N704), .A1(n971), .B0(N692), .B1(n972), .Y(n995) );
  OAI211X1 U1200 ( .A0(n997), .A1(n998), .B0(n953), .C0(n999), .Y(n996) );
  NAND2X1 U1201 ( .A(N745), .B(n973), .Y(n994) );
  OR4X1 U1202 ( .A(n107), .B(n108), .C(n106), .D(n1001), .Y(n997) );
  OR4X1 U1203 ( .A(n112), .B(n111), .C(n110), .D(n109), .Y(n1001) );
  NAND2BX1 U1204 ( .AN(n951), .B(n953), .Y(n948) );
  NAND2X1 U1205 ( .A(n998), .B(n1004), .Y(n951) );
  OAI21XL U1206 ( .A0(n808), .A1(n903), .B0(n1005), .Y(n1004) );
  OAI21XL U1207 ( .A0(n1033), .A1(n1006), .B0(n1007), .Y(n395) );
  NAND2X1 U1208 ( .A(n1008), .B(n1007), .Y(n394) );
  CLKINVX1 U1209 ( .A(n832), .Y(n952) );
  NOR3X1 U1210 ( .A(n833), .B(n1002), .C(n1009), .Y(n832) );
  NOR2X1 U1211 ( .A(n1009), .B(n1002), .Y(n1010) );
  NOR2X1 U1212 ( .A(n785), .B(n800), .Y(n1009) );
  CLKINVX1 U1213 ( .A(n787), .Y(n800) );
  NAND4X1 U1214 ( .A(n68), .B(n55), .C(n959), .D(n778), .Y(n787) );
  NAND4X1 U1215 ( .A(N154), .B(N153), .C(N155), .D(n1012), .Y(n961) );
  NOR3X1 U1216 ( .A(n79), .B(n81), .C(n80), .Y(n1012) );
  NOR4X1 U1217 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(n959) );
  NAND2X1 U1218 ( .A(n1013), .B(n1007), .Y(n392) );
  NAND2X1 U1219 ( .A(n1000), .B(n1006), .Y(n1007) );
  NAND2X1 U1220 ( .A(n1011), .B(n1014), .Y(n1006) );
  OAI21XL U1221 ( .A0(n833), .A1(n801), .B0(n1106), .Y(n1014) );
  CLKINVX1 U1222 ( .A(n831), .Y(n801) );
  NAND2X1 U1223 ( .A(n1003), .B(n903), .Y(n831) );
  CLKINVX1 U1224 ( .A(n999), .Y(n903) );
  NAND2X1 U1225 ( .A(state[0]), .B(n1015), .Y(n999) );
  OAI31XL U1226 ( .A0(n1000), .A1(n1002), .A2(n830), .B0(n1106), .Y(n1011) );
  CLKINVX1 U1227 ( .A(n785), .Y(n830) );
  NAND2X1 U1228 ( .A(n1005), .B(n806), .Y(n785) );
  NOR2X1 U1229 ( .A(n1015), .B(n783), .Y(n806) );
  AND2X1 U1230 ( .A(n955), .B(n1003), .Y(n1002) );
  CLKINVX1 U1231 ( .A(n998), .Y(n1000) );
  NAND2X1 U1232 ( .A(n955), .B(n1005), .Y(n998) );
  NOR3X1 U1233 ( .A(state[2]), .B(state[3]), .C(n788), .Y(n1005) );
  NOR2X1 U1234 ( .A(n1015), .B(state[0]), .Y(n955) );
  AND2X1 U1235 ( .A(n808), .B(n1003), .Y(n833) );
  NOR3X1 U1236 ( .A(n799), .B(state[4]), .C(n797), .Y(n1003) );
endmodule

